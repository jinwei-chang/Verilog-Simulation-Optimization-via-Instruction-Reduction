module dut (out, in);
	output[29:0] out;
	input[49:0] in;
	wire xformtmp6;
	assign xformtmp6 = in[14] ^ in[27];
	wire xformtmp2;
	assign xformtmp2 = in[32] ^ ~xformtmp6;
	wire xformtmp1;
	assign xformtmp1 = xformtmp2 | ~in[14];
	wire xformtmp3;
	assign xformtmp3 = in[20] | in[7];
	assign out[0] = ~xformtmp1 ^ xformtmp3;
	wire xformtmp45;
	assign xformtmp45 = in[33] ^ in[47];
	wire xformtmp52;
	assign xformtmp52 = xformtmp45 | in[49];
	wire xformtmp40;
	assign xformtmp40 = in[39] | in[35];
	wire xformtmp37;
	assign xformtmp37 = in[34] ^ in[35];
	wire xformtmp18;
	assign xformtmp18 = in[45] ^ xformtmp37;
	wire xformtmp38;
	assign xformtmp38 = xformtmp18 & in[13];
	wire xformtmp10;
	assign xformtmp10 = xformtmp40 ^ xformtmp38;
	wire xformtmp17;
	assign xformtmp17 = xformtmp52 & xformtmp10;
	wire xformtmp29;
	assign xformtmp29 = in[19] & in[10];
	wire xformtmp11;
	assign xformtmp11 = xformtmp29 & in[15];
	wire xformtmp14;
	assign xformtmp14 = in[22] & in[25];
	wire xformtmp16;
	assign xformtmp16 = in[24] | in[46];
	wire xformtmp13;
	assign xformtmp13 = xformtmp14 | xformtmp16;
	wire xformtmp8;
	assign xformtmp8 = xformtmp11 & xformtmp13;
	wire xformtmp46;
	assign xformtmp46 = in[1] ^ in[48];
	wire xformtmp44;
	assign xformtmp44 = in[40] | xformtmp46;
	wire xformtmp49;
	assign xformtmp49 = xformtmp8 & xformtmp44;
	wire xformtmp23;
	assign xformtmp23 = in[22] ^ in[5];
	wire xformtmp15;
	assign xformtmp15 = in[18] ^ xformtmp23;
	wire xformtmp9;
	assign xformtmp9 = in[42] | xformtmp15;
	wire xformtmp25;
	assign xformtmp25 = in[16] | xformtmp9;
	wire xformtmp31;
	assign xformtmp31 = xformtmp25 | in[6];
	wire xformtmp27;
	assign xformtmp27 = in[42] & in[12];
	wire xformtmp48;
	assign xformtmp48 = xformtmp31 | xformtmp27;
	wire xformtmp47;
	assign xformtmp47 = in[28] & in[31];
	wire xformtmp30;
	assign xformtmp30 = xformtmp48 | ~xformtmp47;
	wire xformtmp34;
	assign xformtmp34 = xformtmp30 & in[16];
	wire xformtmp35;
	assign xformtmp35 = in[0] | xformtmp34;
	wire xformtmp39;
	assign xformtmp39 = in[28] ^ xformtmp35;
	wire xformtmp36;
	assign xformtmp36 = in[17] | in[39];
	wire xformtmp33;
	assign xformtmp33 = in[38] | xformtmp36;
	wire xformtmp26;
	assign xformtmp26 = xformtmp33 & in[11];
	wire xformtmp22;
	assign xformtmp22 = in[29] & in[9];
	wire xformtmp41;
	assign xformtmp41 = xformtmp26 | xformtmp22;
	wire xformtmp28;
	assign xformtmp28 = xformtmp41 & in[48];
	wire xformtmp19;
	assign xformtmp19 = in[34] ^ in[33];
	wire xformtmp24;
	assign xformtmp24 = xformtmp19 | in[11];
	wire xformtmp43;
	assign xformtmp43 = xformtmp24 & in[44];
	wire xformtmp42;
	assign xformtmp42 = xformtmp43 ^ in[37];
	wire xformtmp50;
	assign xformtmp50 = xformtmp28 | xformtmp42;
	wire xformtmp21;
	assign xformtmp21 = xformtmp39 & xformtmp50;
	wire xformtmp51;
	assign xformtmp51 = xformtmp49 & xformtmp21;
	wire xformtmp12;
	assign xformtmp12 = xformtmp51 | in[5];
	assign out[1] = xformtmp17 & xformtmp12;
	wire xformtmp54;
	assign xformtmp54 = in[41] ^ in[21];
	wire xformtmp58;
	assign xformtmp58 = in[36] ^ xformtmp54;
	wire xformtmp59;
	assign xformtmp59 = in[26] ^ in[23];
	wire xformtmp57;
	assign xformtmp57 = xformtmp59 | in[30];
	wire xformtmp53;
	assign xformtmp53 = in[41] & in[43];
	wire xformtmp55;
	assign xformtmp55 = in[4] & in[8];
	wire xformtmp60;
	assign xformtmp60 = xformtmp53 & xformtmp55;
	wire xformtmp56;
	assign xformtmp56 = xformtmp57 | xformtmp60;
	assign out[2] = xformtmp58 & xformtmp56;
	assign out[3] = ~in[3];
	assign out[4] = 1'b1;
	assign out[5] = 1'b0;
	assign out[6] = 1'b1;
	assign out[7] = 1'b0;
	assign out[8] = 1'b0;
	assign out[9] = 1'b1;
	assign out[10] = 1'b0;
	assign out[11] = 1'b1;
	assign out[12] = 1'b1;
	assign out[13] = 1'b1;
	assign out[14] = 1'b0;
	assign out[15] = 1'b1;
	assign out[16] = 1'b0;
	assign out[17] = 1'b0;
	assign out[18] = 1'b1;
	assign out[19] = 1'b0;
	assign out[20] = 1'b1;
	assign out[21] = 1'b0;
	assign out[22] = 1'b1;
	assign out[23] = 1'b0;
	assign out[24] = 1'b1;
	assign out[25] = 1'b0;
	assign out[26] = 1'b1;
	assign out[27] = 1'b0;
	assign out[28] = 1'b0;
	assign out[29] = 1'b1 ^ in[2];
endmodule

module tb();
    reg[29:0] results[1];
    reg[49:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%50b]", data[0]);
        #1
        $display("results = [%30b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
