module dut (out, in);
	output[29:0] out;
	input[49:0] in;
	wire xformtmp6;
	assign xformtmp6 = in[14] ^ in[27];
	wire xformtmp4;
	assign xformtmp4 = ~xformtmp6;
	wire xformtmp2;
	assign xformtmp2 = in[32] ^ xformtmp4;
	wire xformtmp5;
	assign xformtmp5 = ~in[14];
	wire xformtmp1;
	assign xformtmp1 = xformtmp2 | xformtmp5;
	wire xformtmp7;
	assign xformtmp7 = ~xformtmp1;
	wire xformtmp3;
	assign xformtmp3 = in[7] | in[20];
	assign out[0] = xformtmp7 ^ xformtmp3;
	wire xformtmp45;
	assign xformtmp45 = in[33] ^ in[47];
	wire xformtmp52;
	assign xformtmp52 = in[49] | xformtmp45;
	wire xformtmp40;
	assign xformtmp40 = in[35] | in[39];
	wire xformtmp37;
	assign xformtmp37 = in[34] ^ in[35];
	wire xformtmp18;
	assign xformtmp18 = in[45] ^ xformtmp37;
	wire xformtmp38;
	assign xformtmp38 = in[13] & xformtmp18;
	wire xformtmp10;
	assign xformtmp10 = xformtmp40 ^ xformtmp38;
	wire xformtmp17;
	assign xformtmp17 = xformtmp52 & xformtmp10;
	wire xformtmp29;
	assign xformtmp29 = in[10] & in[19];
	wire xformtmp11;
	assign xformtmp11 = in[15] & xformtmp29;
	wire xformtmp14;
	assign xformtmp14 = in[22] & in[25];
	wire xformtmp16;
	assign xformtmp16 = in[24] | in[46];
	wire xformtmp13;
	assign xformtmp13 = xformtmp14 | xformtmp16;
	wire xformtmp8;
	assign xformtmp8 = xformtmp11 & xformtmp13;
	wire xformtmp46;
	assign xformtmp46 = in[1] ^ in[48];
	wire xformtmp44;
	assign xformtmp44 = in[40] | xformtmp46;
	wire xformtmp49;
	assign xformtmp49 = xformtmp8 & xformtmp44;
	wire xformtmp23;
	assign xformtmp23 = in[5] ^ in[22];
	wire xformtmp15;
	assign xformtmp15 = in[18] ^ xformtmp23;
	wire xformtmp9;
	assign xformtmp9 = in[42] | xformtmp15;
	wire xformtmp25;
	assign xformtmp25 = in[16] | xformtmp9;
	wire xformtmp31;
	assign xformtmp31 = in[6] | xformtmp25;
	wire xformtmp27;
	assign xformtmp27 = in[12] & in[42];
	wire xformtmp48;
	assign xformtmp48 = xformtmp31 | xformtmp27;
	wire xformtmp47;
	assign xformtmp47 = in[28] & in[31];
	wire xformtmp20;
	assign xformtmp20 = ~xformtmp47;
	wire xformtmp30;
	assign xformtmp30 = xformtmp48 | xformtmp20;
	wire xformtmp34;
	assign xformtmp34 = in[16] & xformtmp30;
	wire xformtmp35;
	assign xformtmp35 = in[0] | xformtmp34;
	wire xformtmp39;
	assign xformtmp39 = in[28] ^ xformtmp35;
	wire xformtmp36;
	assign xformtmp36 = in[17] | in[39];
	wire xformtmp33;
	assign xformtmp33 = in[38] | xformtmp36;
	wire xformtmp26;
	assign xformtmp26 = in[11] & xformtmp33;
	wire xformtmp22;
	assign xformtmp22 = in[9] & in[29];
	wire xformtmp41;
	assign xformtmp41 = xformtmp26 | xformtmp22;
	wire xformtmp28;
	assign xformtmp28 = in[48] & xformtmp41;
	wire xformtmp19;
	assign xformtmp19 = in[33] ^ in[34];
	wire xformtmp24;
	assign xformtmp24 = in[11] | xformtmp19;
	wire xformtmp43;
	assign xformtmp43 = in[44] & xformtmp24;
	wire xformtmp42;
	assign xformtmp42 = in[37] ^ xformtmp43;
	wire xformtmp50;
	assign xformtmp50 = xformtmp28 | xformtmp42;
	wire xformtmp21;
	assign xformtmp21 = xformtmp39 & xformtmp50;
	wire xformtmp51;
	assign xformtmp51 = xformtmp49 & xformtmp21;
	wire xformtmp12;
	assign xformtmp12 = in[5] | xformtmp51;
	assign out[1] = xformtmp17 & xformtmp12;
	wire xformtmp54;
	assign xformtmp54 = in[21] ^ in[41];
	wire xformtmp58;
	assign xformtmp58 = in[36] ^ xformtmp54;
	wire xformtmp59;
	assign xformtmp59 = in[23] ^ in[26];
	wire xformtmp57;
	assign xformtmp57 = in[30] | xformtmp59;
	wire xformtmp53;
	assign xformtmp53 = in[41] & in[43];
	wire xformtmp55;
	assign xformtmp55 = in[4] & in[8];
	wire xformtmp60;
	assign xformtmp60 = xformtmp53 & xformtmp55;
	wire xformtmp56;
	assign xformtmp56 = xformtmp57 | xformtmp60;
	assign out[2] = xformtmp58 & xformtmp56;
	assign out[3] = ~in[3];
	assign out[26:4] = 23'b10101010100101110100101;
	wire xformtmp70;
	assign xformtmp70 = 2'b00;
	assign out[28:27] = xformtmp70;
	assign out[29] = ~in[2];
endmodule

module tb();
    reg[29:0] results[1];
    reg[49:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%50b]", data[0]);
        #1
        $display("results = [%30b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
