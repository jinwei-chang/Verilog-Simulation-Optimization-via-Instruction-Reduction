module dut (out, in);
	output[499:0] out;
	input[1499:0] in;
	wire origtmp1;
	wire origtmp2;
	wire origtmp3;
	wire origtmp4;
	wire origtmp5;
	wire origtmp6;
	wire origtmp7;
	wire origtmp8;
	wire origtmp9;
	wire origtmp10;
	wire origtmp11;
	wire origtmp12;
	wire origtmp13;
	wire origtmp14;
	wire origtmp15;
	wire origtmp16;
	wire origtmp17;
	wire origtmp18;
	wire origtmp19;
	wire origtmp20;
	wire origtmp21;
	wire origtmp22;
	wire origtmp23;
	wire origtmp24;
	wire origtmp25;
	wire origtmp26;
	wire origtmp27;
	wire origtmp28;
	wire origtmp29;
	wire origtmp30;
	wire origtmp31;
	wire origtmp32;
	wire origtmp33;
	wire origtmp34;
	wire origtmp35;
	wire origtmp36;
	wire origtmp37;
	wire origtmp38;
	wire origtmp39;
	wire origtmp40;
	wire origtmp41;
	wire origtmp42;
	wire origtmp43;
	wire origtmp44;
	wire origtmp45;
	wire origtmp46;
	wire origtmp47;
	wire origtmp48;
	wire origtmp49;
	wire origtmp50;
	wire origtmp51;
	wire origtmp52;
	wire origtmp53;
	wire origtmp54;
	wire origtmp55;
	wire origtmp56;
	wire origtmp57;
	wire origtmp58;
	wire origtmp59;
	wire origtmp60;
	wire origtmp61;
	wire origtmp62;
	wire origtmp63;
	wire origtmp64;
	wire origtmp65;
	wire origtmp66;
	wire origtmp67;
	wire origtmp68;
	wire origtmp69;
	wire origtmp70;
	wire origtmp71;
	wire origtmp72;
	wire origtmp73;
	wire origtmp74;
	wire origtmp75;
	wire origtmp76;
	wire origtmp77;
	wire origtmp78;
	wire origtmp79;
	wire origtmp80;
	wire origtmp81;
	wire origtmp82;
	wire origtmp83;
	wire origtmp84;
	wire origtmp85;
	wire origtmp86;
	wire origtmp87;
	wire origtmp88;
	wire origtmp89;
	wire origtmp90;
	wire origtmp91;
	wire origtmp92;
	wire origtmp93;
	wire origtmp94;
	wire origtmp95;
	wire origtmp96;
	wire origtmp97;
	wire origtmp98;
	wire origtmp99;
	wire origtmp100;
	wire origtmp101;
	wire origtmp102;
	wire origtmp103;
	wire origtmp104;
	wire origtmp105;
	wire origtmp106;
	wire origtmp107;
	wire origtmp108;
	wire origtmp109;
	wire origtmp110;
	wire origtmp111;
	wire origtmp112;
	wire origtmp113;
	wire origtmp114;
	wire origtmp115;
	wire origtmp116;
	wire origtmp117;
	wire origtmp118;
	wire origtmp119;
	wire origtmp120;
	wire origtmp121;
	wire origtmp122;
	wire origtmp123;
	wire origtmp124;
	wire origtmp125;
	wire origtmp126;
	wire origtmp127;
	wire origtmp128;
	wire origtmp129;
	wire origtmp130;
	wire origtmp131;
	wire origtmp132;
	wire origtmp133;
	wire origtmp134;
	wire origtmp135;
	wire origtmp136;
	wire origtmp137;
	wire origtmp138;
	wire origtmp139;
	wire origtmp140;
	wire origtmp141;
	wire origtmp142;
	wire origtmp143;
	wire origtmp144;
	wire origtmp145;
	wire origtmp146;
	wire origtmp147;
	wire origtmp148;
	wire origtmp149;
	wire origtmp150;
	wire origtmp151;
	wire origtmp152;
	wire origtmp153;
	wire origtmp154;
	wire origtmp155;
	wire origtmp156;
	wire origtmp157;
	wire origtmp158;
	wire origtmp159;
	wire origtmp160;
	wire origtmp161;
	wire origtmp162;
	wire origtmp163;
	wire origtmp164;
	wire origtmp165;
	wire origtmp166;
	wire origtmp167;
	wire origtmp168;
	wire origtmp169;
	wire origtmp170;
	wire origtmp171;
	wire origtmp172;
	wire origtmp173;
	wire origtmp174;
	wire origtmp175;
	wire origtmp176;
	wire origtmp177;
	wire origtmp178;
	wire origtmp179;
	wire origtmp180;
	wire origtmp181;
	wire origtmp182;
	wire origtmp183;
	wire origtmp184;
	wire origtmp185;
	wire origtmp186;
	wire origtmp187;
	wire origtmp188;
	wire origtmp189;
	wire origtmp190;
	wire origtmp191;
	wire origtmp192;
	wire origtmp193;
	wire origtmp194;
	wire origtmp195;
	wire origtmp196;
	wire origtmp197;
	wire origtmp198;
	wire origtmp199;
	wire origtmp200;
	wire origtmp201;
	wire origtmp202;
	wire origtmp203;
	wire origtmp204;
	wire origtmp205;
	wire origtmp206;
	wire origtmp207;
	wire origtmp208;
	wire origtmp209;
	wire origtmp210;
	wire origtmp211;
	wire origtmp212;
	wire origtmp213;
	wire origtmp214;
	wire origtmp215;
	wire origtmp216;
	wire origtmp217;
	wire origtmp218;
	wire origtmp219;
	wire origtmp220;
	wire origtmp221;
	wire origtmp222;
	wire origtmp223;
	wire origtmp224;
	wire origtmp225;
	wire origtmp226;
	wire origtmp227;
	wire origtmp228;
	wire origtmp229;
	wire origtmp230;
	wire origtmp231;
	wire origtmp232;
	wire origtmp233;
	wire origtmp234;
	wire origtmp235;
	wire origtmp236;
	wire origtmp237;
	wire origtmp238;
	wire origtmp239;
	wire origtmp240;
	wire origtmp241;
	wire origtmp242;
	wire origtmp243;
	wire origtmp244;
	wire origtmp245;
	wire origtmp246;
	wire origtmp247;
	wire origtmp248;
	wire origtmp249;
	wire origtmp250;
	wire origtmp251;
	wire origtmp252;
	wire origtmp253;
	wire origtmp254;
	wire origtmp255;
	wire origtmp256;
	wire origtmp257;
	wire origtmp258;
	wire origtmp259;
	wire origtmp260;
	wire origtmp261;
	wire origtmp262;
	wire origtmp263;
	wire origtmp264;
	wire origtmp265;
	wire origtmp266;
	wire origtmp267;
	wire origtmp268;
	wire origtmp269;
	wire origtmp270;
	wire origtmp271;
	wire origtmp272;
	wire origtmp273;
	wire origtmp274;
	wire origtmp275;
	wire origtmp276;
	wire origtmp277;
	wire origtmp278;
	wire origtmp279;
	wire origtmp280;
	wire origtmp281;
	wire origtmp282;
	wire origtmp283;
	wire origtmp284;
	wire origtmp285;
	wire origtmp286;
	wire origtmp287;
	wire origtmp288;
	wire origtmp289;
	wire origtmp290;
	wire origtmp291;
	wire origtmp292;
	wire origtmp293;
	wire origtmp294;
	wire origtmp295;
	wire origtmp296;
	wire origtmp297;
	wire origtmp298;
	wire origtmp299;
	wire origtmp300;
	wire origtmp301;
	wire origtmp302;
	wire origtmp303;
	wire origtmp304;
	wire origtmp305;
	wire origtmp306;
	wire origtmp307;
	wire origtmp308;
	wire origtmp309;
	wire origtmp310;
	wire origtmp311;
	wire origtmp312;
	wire origtmp313;
	wire origtmp314;
	wire origtmp315;
	wire origtmp316;
	wire origtmp317;
	wire origtmp318;
	wire origtmp319;
	wire origtmp320;
	wire origtmp321;
	wire origtmp322;
	wire origtmp323;
	wire origtmp324;
	wire origtmp325;
	wire origtmp326;
	wire origtmp327;
	wire origtmp328;
	wire origtmp329;
	wire origtmp330;
	wire origtmp331;
	wire origtmp332;
	wire origtmp333;
	wire origtmp334;
	wire origtmp335;
	wire origtmp336;
	wire origtmp337;
	wire origtmp338;
	wire origtmp339;
	wire origtmp340;
	wire origtmp341;
	wire origtmp342;
	wire origtmp343;
	wire origtmp344;
	wire origtmp345;
	wire origtmp346;
	wire origtmp347;
	wire origtmp348;
	wire origtmp349;
	wire origtmp350;
	wire origtmp351;
	wire origtmp352;
	wire origtmp353;
	wire origtmp354;
	wire origtmp355;
	wire origtmp356;
	wire origtmp357;
	wire origtmp358;
	wire origtmp359;
	wire origtmp360;
	wire origtmp361;
	wire origtmp362;
	wire origtmp363;
	wire origtmp364;
	wire origtmp365;
	wire origtmp366;
	wire origtmp367;
	wire origtmp368;
	wire origtmp369;
	wire origtmp370;
	wire origtmp371;
	wire origtmp372;
	wire origtmp373;
	wire origtmp374;
	wire origtmp375;
	wire origtmp376;
	wire origtmp377;
	wire origtmp378;
	wire origtmp379;
	wire origtmp380;
	wire origtmp381;
	wire origtmp382;
	wire origtmp383;
	wire origtmp384;
	wire origtmp385;
	wire origtmp386;
	wire origtmp387;
	wire origtmp388;
	wire origtmp389;
	wire origtmp390;
	wire origtmp391;
	wire origtmp392;
	wire origtmp393;
	wire origtmp394;
	wire origtmp395;
	wire origtmp396;
	wire origtmp397;
	wire origtmp398;
	wire origtmp399;
	wire origtmp400;
	wire origtmp401;
	wire origtmp402;
	wire origtmp403;
	wire origtmp404;
	wire origtmp405;
	wire origtmp406;
	wire origtmp407;
	wire origtmp408;
	wire origtmp409;
	wire origtmp410;
	wire origtmp411;
	wire origtmp412;
	wire origtmp413;
	wire origtmp414;
	wire origtmp415;
	wire origtmp416;
	wire origtmp417;
	wire origtmp418;
	wire origtmp419;
	wire origtmp420;
	wire origtmp421;
	wire origtmp422;
	wire origtmp423;
	wire origtmp424;
	wire origtmp425;
	wire origtmp426;
	wire origtmp427;
	wire origtmp428;
	wire origtmp429;
	wire origtmp430;
	wire origtmp431;
	wire origtmp432;
	wire origtmp433;
	wire origtmp434;
	wire origtmp435;
	wire origtmp436;
	wire origtmp437;
	wire origtmp438;
	wire origtmp439;
	wire origtmp440;
	wire origtmp441;
	wire origtmp442;
	wire origtmp443;
	wire origtmp444;
	wire origtmp445;
	wire origtmp446;
	wire origtmp447;
	wire origtmp448;
	wire origtmp449;
	wire origtmp450;
	wire origtmp451;
	wire origtmp452;
	wire origtmp453;
	wire origtmp454;
	wire origtmp455;
	wire origtmp456;
	wire origtmp457;
	wire origtmp458;
	wire origtmp459;
	wire origtmp460;
	wire origtmp461;
	wire origtmp462;
	wire origtmp463;
	wire origtmp464;
	wire origtmp465;
	wire origtmp466;
	wire origtmp467;
	wire origtmp468;
	wire origtmp469;
	wire origtmp470;
	wire origtmp471;
	wire origtmp472;
	wire origtmp473;
	wire origtmp474;
	wire origtmp475;
	wire origtmp476;
	wire origtmp477;
	wire origtmp478;
	wire origtmp479;
	wire origtmp480;
	wire origtmp481;
	wire origtmp482;
	wire origtmp483;
	wire origtmp484;
	wire origtmp485;
	wire origtmp486;
	wire origtmp487;
	wire origtmp488;
	wire origtmp489;
	wire origtmp490;
	wire origtmp491;
	wire origtmp492;
	wire origtmp493;
	wire origtmp494;
	wire origtmp495;
	wire origtmp496;
	wire origtmp497;
	wire origtmp498;
	wire origtmp499;
	wire origtmp500;
	wire origtmp501;
	wire origtmp502;
	wire origtmp503;
	wire origtmp504;
	wire origtmp505;
	wire origtmp506;
	wire origtmp507;
	wire origtmp508;
	wire origtmp509;
	wire origtmp510;
	wire origtmp511;
	wire origtmp512;
	wire origtmp513;
	wire origtmp514;
	wire origtmp515;
	wire origtmp516;
	wire origtmp517;
	wire origtmp518;
	wire origtmp519;
	wire origtmp520;
	wire origtmp521;
	wire origtmp522;
	wire origtmp523;
	wire origtmp524;
	wire origtmp525;
	wire origtmp526;
	wire origtmp527;
	wire origtmp528;
	wire origtmp529;
	wire origtmp530;
	wire origtmp531;
	wire origtmp532;
	wire origtmp533;
	wire origtmp534;
	wire origtmp535;
	wire origtmp536;
	wire origtmp537;
	wire origtmp538;
	wire origtmp539;
	wire origtmp540;
	wire origtmp541;
	wire origtmp542;
	wire origtmp543;
	wire origtmp544;
	wire origtmp545;
	wire origtmp546;
	wire origtmp547;
	wire origtmp548;
	wire origtmp549;
	wire origtmp550;
	wire origtmp551;
	wire origtmp552;
	wire origtmp553;
	wire origtmp554;
	wire origtmp555;
	wire origtmp556;
	wire origtmp557;
	wire origtmp558;
	wire origtmp559;
	wire origtmp560;
	wire origtmp561;
	wire origtmp562;
	wire origtmp563;
	wire origtmp564;
	wire origtmp565;
	wire origtmp566;
	wire origtmp567;
	wire origtmp568;
	wire origtmp569;
	wire origtmp570;
	wire origtmp571;
	wire origtmp572;
	wire origtmp573;
	wire origtmp574;
	wire origtmp575;
	wire origtmp576;
	wire origtmp577;
	wire origtmp578;
	wire origtmp579;
	wire origtmp580;
	wire origtmp581;
	wire origtmp582;
	wire origtmp583;
	wire origtmp584;
	wire origtmp585;
	wire origtmp586;
	wire origtmp587;
	wire origtmp588;
	wire origtmp589;
	wire origtmp590;
	wire origtmp591;
	wire origtmp592;
	wire origtmp593;
	wire origtmp594;
	wire origtmp595;
	wire origtmp596;
	wire origtmp597;
	wire origtmp598;
	wire origtmp599;
	wire origtmp600;
	wire origtmp601;
	wire origtmp602;
	wire origtmp603;
	wire origtmp604;
	wire origtmp605;
	wire origtmp606;
	wire origtmp607;
	wire origtmp608;
	wire origtmp609;
	wire origtmp610;
	wire origtmp611;
	wire origtmp612;
	wire origtmp613;
	wire origtmp614;
	wire origtmp615;
	wire origtmp616;
	wire origtmp617;
	wire origtmp618;
	wire origtmp619;
	wire origtmp620;
	wire origtmp621;
	wire origtmp622;
	wire origtmp623;
	wire origtmp624;
	wire origtmp625;
	wire origtmp626;
	wire origtmp627;
	wire origtmp628;
	wire origtmp629;
	wire origtmp630;
	wire origtmp631;
	wire origtmp632;
	wire origtmp633;
	wire origtmp634;
	wire origtmp635;
	wire origtmp636;
	wire origtmp637;
	wire origtmp638;
	wire origtmp639;
	wire origtmp640;
	wire origtmp641;
	wire origtmp642;
	wire origtmp643;
	wire origtmp644;
	wire origtmp645;
	wire origtmp646;
	wire origtmp647;
	wire origtmp648;
	wire origtmp649;
	wire origtmp650;
	wire origtmp651;
	wire origtmp652;
	wire origtmp653;
	wire origtmp654;
	wire origtmp655;
	wire origtmp656;
	wire origtmp657;
	wire origtmp658;
	wire origtmp659;
	wire origtmp660;
	wire origtmp661;
	wire origtmp662;
	wire origtmp663;
	wire origtmp664;
	wire origtmp665;
	wire origtmp666;
	wire origtmp667;
	wire origtmp668;
	wire origtmp669;
	wire origtmp670;
	wire origtmp671;
	wire origtmp672;
	wire origtmp673;
	wire origtmp674;
	wire origtmp675;
	wire origtmp676;
	wire origtmp677;
	wire origtmp678;
	wire origtmp679;
	wire origtmp680;
	wire origtmp681;
	wire origtmp682;
	wire origtmp683;
	wire origtmp684;
	wire origtmp685;
	wire origtmp686;
	wire origtmp687;
	wire origtmp688;
	wire origtmp689;
	wire origtmp690;
	wire origtmp691;
	wire origtmp692;
	wire origtmp693;
	wire origtmp694;
	wire origtmp695;
	wire origtmp696;
	wire origtmp697;
	wire origtmp698;
	wire origtmp699;
	wire origtmp700;
	wire origtmp701;
	wire origtmp702;
	wire origtmp703;
	wire origtmp704;
	wire origtmp705;
	wire origtmp706;
	wire origtmp707;
	wire origtmp708;
	wire origtmp709;
	wire origtmp710;
	wire origtmp711;
	wire origtmp712;
	wire origtmp713;
	wire origtmp714;
	wire origtmp715;
	wire origtmp716;
	wire origtmp717;
	wire origtmp718;
	wire origtmp719;
	wire origtmp720;
	wire origtmp721;
	wire origtmp722;
	wire origtmp723;
	wire origtmp724;
	wire origtmp725;
	wire origtmp726;
	wire origtmp727;
	wire origtmp728;
	wire origtmp729;
	wire origtmp730;
	wire origtmp731;
	wire origtmp732;
	wire origtmp733;
	wire origtmp734;
	wire origtmp735;
	wire origtmp736;
	wire origtmp737;
	wire origtmp738;
	wire origtmp739;
	wire origtmp740;
	wire origtmp741;
	wire origtmp742;
	wire origtmp743;
	wire origtmp744;
	wire origtmp745;
	wire origtmp746;
	wire origtmp747;
	wire origtmp748;
	wire origtmp749;
	wire origtmp750;
	wire origtmp751;
	wire origtmp752;
	wire origtmp753;
	wire origtmp754;
	wire origtmp755;
	wire origtmp756;
	wire origtmp757;
	wire origtmp758;
	wire origtmp759;
	wire origtmp760;
	wire origtmp761;
	wire origtmp762;
	wire origtmp763;
	wire origtmp764;
	wire origtmp765;
	wire origtmp766;
	wire origtmp767;
	wire origtmp768;
	wire origtmp769;
	wire origtmp770;
	wire origtmp771;
	wire origtmp772;
	wire origtmp773;
	wire origtmp774;
	wire origtmp775;
	wire origtmp776;
	wire origtmp777;
	wire origtmp778;
	wire origtmp779;
	wire origtmp780;
	wire origtmp781;
	wire origtmp782;
	wire origtmp783;
	wire origtmp784;
	wire origtmp785;
	wire origtmp786;
	wire origtmp787;
	wire origtmp788;
	wire origtmp789;
	wire origtmp790;
	wire origtmp791;
	wire origtmp792;
	wire origtmp793;
	wire origtmp794;
	wire origtmp795;
	wire origtmp796;
	wire origtmp797;
	wire origtmp798;
	wire origtmp799;
	wire origtmp800;
	wire origtmp801;
	wire origtmp802;
	wire origtmp803;
	wire origtmp804;
	wire origtmp805;
	wire origtmp806;
	wire origtmp807;
	wire origtmp808;
	wire origtmp809;
	wire origtmp810;
	wire origtmp811;
	wire origtmp812;
	wire origtmp813;
	wire origtmp814;
	wire origtmp815;
	wire origtmp816;
	wire origtmp817;
	wire origtmp818;
	wire origtmp819;
	wire origtmp820;
	wire origtmp821;
	wire origtmp822;
	wire origtmp823;
	wire origtmp824;
	wire origtmp825;
	wire origtmp826;
	wire origtmp827;
	wire origtmp828;
	wire origtmp829;
	wire origtmp830;
	wire origtmp831;
	wire origtmp832;
	wire origtmp833;
	wire origtmp834;
	wire origtmp835;
	wire origtmp836;
	wire origtmp837;
	wire origtmp838;
	wire origtmp839;
	wire origtmp840;
	wire origtmp841;
	wire origtmp842;
	wire origtmp843;
	wire origtmp844;
	wire origtmp845;
	wire origtmp846;
	wire origtmp847;
	wire origtmp848;
	wire origtmp849;
	wire origtmp850;
	wire origtmp851;
	wire origtmp852;
	wire origtmp853;
	wire origtmp854;
	wire origtmp855;
	wire origtmp856;
	wire origtmp857;
	wire origtmp858;
	wire origtmp859;
	wire origtmp860;
	wire origtmp861;
	wire origtmp862;
	wire origtmp863;
	wire origtmp864;
	wire origtmp865;
	wire origtmp866;
	wire origtmp867;
	wire origtmp868;
	wire origtmp869;
	wire origtmp870;
	wire origtmp871;
	wire origtmp872;
	wire origtmp873;
	wire origtmp874;
	wire origtmp875;
	wire origtmp876;
	wire origtmp877;
	wire origtmp878;
	wire origtmp879;
	wire origtmp880;
	wire origtmp881;
	wire origtmp882;
	wire origtmp883;
	wire origtmp884;
	wire origtmp885;
	wire origtmp886;
	wire origtmp887;
	wire origtmp888;
	wire origtmp889;
	wire origtmp890;
	wire origtmp891;
	wire origtmp892;
	wire origtmp893;
	wire origtmp894;
	wire origtmp895;
	wire origtmp896;
	wire origtmp897;
	wire origtmp898;
	wire origtmp899;
	wire origtmp900;
	wire origtmp901;
	wire origtmp902;
	wire origtmp903;
	wire origtmp904;
	wire origtmp905;
	wire origtmp906;
	wire origtmp907;
	wire origtmp908;
	wire origtmp909;
	wire origtmp910;
	wire origtmp911;
	wire origtmp912;
	wire origtmp913;
	wire origtmp914;
	wire origtmp915;
	wire origtmp916;
	wire origtmp917;
	wire origtmp918;
	wire origtmp919;
	wire origtmp920;
	wire origtmp921;
	wire origtmp922;
	wire origtmp923;
	wire origtmp924;
	wire origtmp925;
	wire origtmp926;
	wire origtmp927;
	wire origtmp928;
	wire origtmp929;
	wire origtmp930;
	wire origtmp931;
	wire origtmp932;
	wire origtmp933;
	wire origtmp934;
	wire origtmp935;
	wire origtmp936;
	wire origtmp937;
	wire origtmp938;
	wire origtmp939;
	wire origtmp940;
	wire origtmp941;
	wire origtmp942;
	wire origtmp943;
	wire origtmp944;
	wire origtmp945;
	wire origtmp946;
	wire origtmp947;
	wire origtmp948;
	wire origtmp949;
	wire origtmp950;
	wire origtmp951;
	wire origtmp952;
	wire origtmp953;
	wire origtmp954;
	wire origtmp955;
	wire origtmp956;
	wire origtmp957;
	wire origtmp958;
	wire origtmp959;
	wire origtmp960;
	wire origtmp961;
	wire origtmp962;
	wire origtmp963;
	wire origtmp964;
	wire origtmp965;
	wire origtmp966;
	wire origtmp967;
	wire origtmp968;
	wire origtmp969;
	wire origtmp970;
	wire origtmp971;
	wire origtmp972;
	wire origtmp973;
	wire origtmp974;
	wire origtmp975;
	wire origtmp976;
	wire origtmp977;
	wire origtmp978;
	wire origtmp979;
	wire origtmp980;
	wire origtmp981;
	wire origtmp982;
	wire origtmp983;
	wire origtmp984;
	wire origtmp985;
	wire origtmp986;
	wire origtmp987;
	wire origtmp988;
	wire origtmp989;
	wire origtmp990;
	wire origtmp991;
	wire origtmp992;
	wire origtmp993;
	wire origtmp994;
	wire origtmp995;
	wire origtmp996;
	wire origtmp997;
	wire origtmp998;
	wire origtmp999;
	wire origtmp1000;
	wire origtmp1001;
	wire origtmp1002;
	wire origtmp1003;
	wire origtmp1004;
	wire origtmp1005;
	wire origtmp1006;
	wire origtmp1007;
	wire origtmp1008;
	wire origtmp1009;
	wire origtmp1010;
	wire origtmp1011;
	wire origtmp1012;
	wire origtmp1013;
	wire origtmp1014;
	wire origtmp1015;
	wire origtmp1016;
	wire origtmp1017;
	wire origtmp1018;
	wire origtmp1019;
	wire origtmp1020;
	wire origtmp1021;
	wire origtmp1022;
	wire origtmp1023;
	wire origtmp1024;
	wire origtmp1025;
	wire origtmp1026;
	wire origtmp1027;
	wire origtmp1028;
	wire origtmp1029;
	wire origtmp1030;
	wire origtmp1031;
	wire origtmp1032;
	wire origtmp1033;
	wire origtmp1034;
	wire origtmp1035;
	wire origtmp1036;
	wire origtmp1037;
	wire origtmp1038;
	wire origtmp1039;
	wire origtmp1040;
	wire origtmp1041;
	wire origtmp1042;
	wire origtmp1043;
	wire origtmp1044;
	wire origtmp1045;
	wire origtmp1046;
	wire origtmp1047;
	wire origtmp1048;
	wire origtmp1049;
	wire origtmp1050;
	wire origtmp1051;
	wire origtmp1052;
	wire origtmp1053;
	wire origtmp1054;
	wire origtmp1055;
	wire origtmp1056;
	wire origtmp1057;
	wire origtmp1058;
	wire origtmp1059;
	wire origtmp1060;
	wire origtmp1061;
	wire origtmp1062;
	wire origtmp1063;
	wire origtmp1064;
	wire origtmp1065;
	wire origtmp1066;
	wire origtmp1067;
	wire origtmp1068;
	wire origtmp1069;
	wire origtmp1070;
	wire origtmp1071;
	wire origtmp1072;
	wire origtmp1073;
	wire origtmp1074;
	wire origtmp1075;
	wire origtmp1076;
	wire origtmp1077;
	wire origtmp1078;
	wire origtmp1079;
	wire origtmp1080;
	wire origtmp1081;
	wire origtmp1082;
	wire origtmp1083;
	wire origtmp1084;
	wire origtmp1085;
	wire origtmp1086;
	wire origtmp1087;
	wire origtmp1088;
	wire origtmp1089;
	wire origtmp1090;
	wire origtmp1091;
	wire origtmp1092;
	wire origtmp1093;
	wire origtmp1094;
	wire origtmp1095;
	wire origtmp1096;
	wire origtmp1097;
	wire origtmp1098;
	wire origtmp1099;
	wire origtmp1100;
	wire origtmp1101;
	wire origtmp1102;
	wire origtmp1103;
	wire origtmp1104;
	wire origtmp1105;
	wire origtmp1106;
	wire origtmp1107;
	wire origtmp1108;
	wire origtmp1109;
	wire origtmp1110;
	wire origtmp1111;
	wire origtmp1112;
	wire origtmp1113;
	wire origtmp1114;
	wire origtmp1115;
	wire origtmp1116;
	wire origtmp1117;
	wire origtmp1118;
	wire origtmp1119;
	wire origtmp1120;
	wire origtmp1121;
	wire origtmp1122;
	wire origtmp1123;
	wire origtmp1124;
	wire origtmp1125;
	wire origtmp1126;
	wire origtmp1127;
	wire origtmp1128;
	wire origtmp1129;
	wire origtmp1130;
	wire origtmp1131;
	wire origtmp1132;
	wire origtmp1133;
	wire origtmp1134;
	wire origtmp1135;
	wire origtmp1136;
	wire origtmp1137;
	wire origtmp1138;
	wire origtmp1139;
	wire origtmp1140;
	wire origtmp1141;
	wire origtmp1142;
	wire origtmp1143;
	wire origtmp1144;
	wire origtmp1145;
	wire origtmp1146;
	wire origtmp1147;
	wire origtmp1148;
	wire origtmp1149;
	wire origtmp1150;
	wire origtmp1151;
	wire origtmp1152;
	wire origtmp1153;
	wire origtmp1154;
	wire origtmp1155;
	wire origtmp1156;
	wire origtmp1157;
	wire origtmp1158;
	wire origtmp1159;
	wire origtmp1160;
	wire origtmp1161;
	wire origtmp1162;
	wire origtmp1163;
	wire origtmp1164;
	wire origtmp1165;
	wire origtmp1166;
	wire origtmp1167;
	wire origtmp1168;
	wire origtmp1169;
	wire origtmp1170;
	wire origtmp1171;
	wire origtmp1172;
	wire origtmp1173;
	wire origtmp1174;
	wire origtmp1175;
	wire origtmp1176;
	wire origtmp1177;
	wire origtmp1178;
	wire origtmp1179;
	wire origtmp1180;
	wire origtmp1181;
	wire origtmp1182;
	wire origtmp1183;
	wire origtmp1184;
	wire origtmp1185;
	wire origtmp1186;
	wire origtmp1187;
	wire origtmp1188;
	wire origtmp1189;
	wire origtmp1190;
	wire origtmp1191;
	wire origtmp1192;
	wire origtmp1193;
	wire origtmp1194;
	wire origtmp1195;
	wire origtmp1196;
	wire origtmp1197;
	wire origtmp1198;
	wire origtmp1199;
	wire origtmp1200;
	wire origtmp1201;
	wire origtmp1202;
	wire origtmp1203;
	wire origtmp1204;
	wire origtmp1205;
	wire origtmp1206;
	wire origtmp1207;
	wire origtmp1208;
	wire origtmp1209;
	wire origtmp1210;
	wire origtmp1211;
	wire origtmp1212;
	wire origtmp1213;
	wire origtmp1214;
	wire origtmp1215;
	wire origtmp1216;
	wire origtmp1217;
	wire origtmp1218;
	wire origtmp1219;
	wire origtmp1220;
	wire origtmp1221;
	wire origtmp1222;
	wire origtmp1223;
	wire origtmp1224;
	wire origtmp1225;
	wire origtmp1226;
	wire origtmp1227;
	wire origtmp1228;
	wire origtmp1229;
	wire origtmp1230;
	wire origtmp1231;
	wire origtmp1232;
	wire origtmp1233;
	wire origtmp1234;
	wire origtmp1235;
	wire origtmp1236;
	wire origtmp1237;
	wire origtmp1238;
	wire origtmp1239;
	wire origtmp1240;
	wire origtmp1241;
	wire origtmp1242;
	wire origtmp1243;
	wire origtmp1244;
	wire origtmp1245;
	wire origtmp1246;
	wire origtmp1247;
	wire origtmp1248;
	wire origtmp1249;
	wire origtmp1250;
	wire origtmp1251;
	wire origtmp1252;
	wire origtmp1253;
	wire origtmp1254;
	wire origtmp1255;
	wire origtmp1256;
	wire origtmp1257;
	wire origtmp1258;
	wire origtmp1259;
	wire origtmp1260;
	wire origtmp1261;
	wire origtmp1262;
	wire origtmp1263;
	wire origtmp1264;
	wire origtmp1265;
	wire origtmp1266;
	wire origtmp1267;
	wire origtmp1268;
	wire origtmp1269;
	wire origtmp1270;
	wire origtmp1271;
	wire origtmp1272;
	wire origtmp1273;
	wire origtmp1274;
	wire origtmp1275;
	wire origtmp1276;
	wire origtmp1277;
	wire origtmp1278;
	wire origtmp1279;
	wire origtmp1280;
	wire origtmp1281;
	wire origtmp1282;
	wire origtmp1283;
	wire origtmp1284;
	wire origtmp1285;
	wire origtmp1286;
	wire origtmp1287;
	wire origtmp1288;
	wire origtmp1289;
	wire origtmp1290;
	wire origtmp1291;
	wire origtmp1292;
	wire origtmp1293;
	wire origtmp1294;
	wire origtmp1295;
	wire origtmp1296;
	wire origtmp1297;
	wire origtmp1298;
	wire origtmp1299;
	wire origtmp1300;
	wire origtmp1301;
	wire origtmp1302;
	wire origtmp1303;
	wire origtmp1304;
	wire origtmp1305;
	wire origtmp1306;
	wire origtmp1307;
	wire origtmp1308;
	wire origtmp1309;
	wire origtmp1310;
	wire origtmp1311;
	wire origtmp1312;
	wire origtmp1313;
	wire origtmp1314;
	wire origtmp1315;
	wire origtmp1316;
	wire origtmp1317;
	wire origtmp1318;
	wire origtmp1319;
	wire origtmp1320;
	wire origtmp1321;
	wire origtmp1322;
	wire origtmp1323;
	wire origtmp1324;
	wire origtmp1325;
	wire origtmp1326;
	wire origtmp1327;
	wire origtmp1328;
	wire origtmp1329;
	wire origtmp1330;
	wire origtmp1331;
	wire origtmp1332;
	wire origtmp1333;
	wire origtmp1334;
	wire origtmp1335;
	wire origtmp1336;
	wire origtmp1337;
	wire origtmp1338;
	wire origtmp1339;
	wire origtmp1340;
	wire origtmp1341;
	wire origtmp1342;
	wire origtmp1343;
	wire origtmp1344;
	wire origtmp1345;
	wire origtmp1346;
	wire origtmp1347;
	wire origtmp1348;
	wire origtmp1349;
	wire origtmp1350;
	wire origtmp1351;
	wire origtmp1352;
	wire origtmp1353;
	wire origtmp1354;
	wire origtmp1355;
	wire origtmp1356;
	wire origtmp1357;
	wire origtmp1358;
	wire origtmp1359;
	wire origtmp1360;
	wire origtmp1361;
	wire origtmp1362;
	wire origtmp1363;
	wire origtmp1364;
	wire origtmp1365;
	wire origtmp1366;
	wire origtmp1367;
	wire origtmp1368;
	wire origtmp1369;
	wire origtmp1370;
	wire origtmp1371;
	wire origtmp1372;
	wire origtmp1373;
	wire origtmp1374;
	wire origtmp1375;
	wire origtmp1376;
	wire origtmp1377;
	wire origtmp1378;
	wire origtmp1379;
	wire origtmp1380;
	wire origtmp1381;
	wire origtmp1382;
	wire origtmp1383;
	wire origtmp1384;
	wire origtmp1385;
	wire origtmp1386;
	wire origtmp1387;
	wire origtmp1388;
	wire origtmp1389;
	wire origtmp1390;
	wire origtmp1391;
	wire origtmp1392;
	wire origtmp1393;
	wire origtmp1394;
	wire origtmp1395;
	wire origtmp1396;
	wire origtmp1397;
	wire origtmp1398;
	wire origtmp1399;
	wire origtmp1400;
	wire origtmp1401;
	wire origtmp1402;
	wire origtmp1403;
	wire origtmp1404;
	wire origtmp1405;
	wire origtmp1406;
	wire origtmp1407;
	wire origtmp1408;
	wire origtmp1409;
	wire origtmp1410;
	wire origtmp1411;
	wire origtmp1412;
	wire origtmp1413;
	wire origtmp1414;
	wire origtmp1415;
	wire origtmp1416;
	wire origtmp1417;
	wire origtmp1418;
	wire origtmp1419;
	wire origtmp1420;
	wire origtmp1421;
	wire origtmp1422;
	wire origtmp1423;
	wire origtmp1424;
	wire origtmp1425;
	wire origtmp1426;
	wire origtmp1427;
	wire origtmp1428;
	wire origtmp1429;
	wire origtmp1430;
	wire origtmp1431;
	wire origtmp1432;
	wire origtmp1433;
	wire origtmp1434;
	wire origtmp1435;
	wire origtmp1436;
	wire origtmp1437;
	wire origtmp1438;
	wire origtmp1439;
	wire origtmp1440;
	wire origtmp1441;
	wire origtmp1442;
	wire origtmp1443;
	wire origtmp1444;
	wire origtmp1445;
	wire origtmp1446;
	wire origtmp1447;
	wire origtmp1448;
	wire origtmp1449;
	wire origtmp1450;
	wire origtmp1451;
	wire origtmp1452;
	wire origtmp1453;
	wire origtmp1454;
	wire origtmp1455;
	wire origtmp1456;
	wire origtmp1457;
	wire origtmp1458;
	wire origtmp1459;
	wire origtmp1460;
	wire origtmp1461;
	wire origtmp1462;
	wire origtmp1463;
	wire origtmp1464;
	wire origtmp1465;
	wire origtmp1466;
	wire origtmp1467;
	wire origtmp1468;
	wire origtmp1469;
	wire origtmp1470;
	wire origtmp1471;
	wire origtmp1472;
	wire origtmp1473;
	wire origtmp1474;
	wire origtmp1475;
	wire origtmp1476;
	wire origtmp1477;
	wire origtmp1478;
	wire origtmp1479;
	wire origtmp1480;
	wire origtmp1481;
	wire origtmp1482;
	wire origtmp1483;
	wire origtmp1484;
	wire origtmp1485;
	wire origtmp1486;
	wire origtmp1487;
	wire origtmp1488;
	wire origtmp1489;
	wire origtmp1490;
	wire origtmp1491;
	wire origtmp1492;
	wire origtmp1493;
	wire origtmp1494;
	wire origtmp1495;
	wire origtmp1496;
	wire origtmp1497;
	wire origtmp1498;
	wire origtmp1499;
	wire origtmp1500;
	wire origtmp1501;
	wire origtmp1502;
	wire origtmp1503;
	wire origtmp1504;
	wire origtmp1505;
	wire origtmp1506;
	wire origtmp1507;
	wire origtmp1508;
	wire origtmp1509;
	wire origtmp1510;
	wire origtmp1511;
	wire origtmp1512;
	wire origtmp1513;
	wire origtmp1514;
	wire origtmp1515;
	wire origtmp1516;
	wire origtmp1517;
	wire origtmp1518;
	wire origtmp1519;
	wire origtmp1520;
	wire origtmp1521;
	wire origtmp1522;
	wire origtmp1523;
	wire origtmp1524;
	wire origtmp1525;
	wire origtmp1526;
	wire origtmp1527;
	wire origtmp1528;
	wire origtmp1529;
	wire origtmp1530;
	wire origtmp1531;
	wire origtmp1532;
	wire origtmp1533;
	wire origtmp1534;
	wire origtmp1535;
	wire origtmp1536;
	wire origtmp1537;
	wire origtmp1538;
	wire origtmp1539;
	wire origtmp1540;
	wire origtmp1541;
	wire origtmp1542;
	wire origtmp1543;
	wire origtmp1544;
	wire origtmp1545;
	wire origtmp1546;
	wire origtmp1547;
	wire origtmp1548;
	wire origtmp1549;
	wire origtmp1550;
	wire origtmp1551;
	wire origtmp1552;
	wire origtmp1553;
	wire origtmp1554;
	wire origtmp1555;
	wire origtmp1556;
	wire origtmp1557;
	wire origtmp1558;
	wire origtmp1559;
	wire origtmp1560;
	wire origtmp1561;
	wire origtmp1562;
	wire origtmp1563;
	wire origtmp1564;
	wire origtmp1565;
	wire origtmp1566;
	wire origtmp1567;
	wire origtmp1568;
	wire origtmp1569;
	wire origtmp1570;
	wire origtmp1571;
	wire origtmp1572;
	wire origtmp1573;
	wire origtmp1574;
	wire origtmp1575;
	wire origtmp1576;
	wire origtmp1577;
	wire origtmp1578;
	wire origtmp1579;
	wire origtmp1580;
	wire origtmp1581;
	wire origtmp1582;
	wire origtmp1583;
	wire origtmp1584;
	wire origtmp1585;
	wire origtmp1586;
	wire origtmp1587;
	wire origtmp1588;
	wire origtmp1589;
	wire origtmp1590;
	wire origtmp1591;
	wire origtmp1592;
	wire origtmp1593;
	wire origtmp1594;
	wire origtmp1595;
	wire origtmp1596;
	wire origtmp1597;
	wire origtmp1598;
	wire origtmp1599;
	wire origtmp1600;
	wire origtmp1601;
	wire origtmp1602;
	wire origtmp1603;
	wire origtmp1604;
	wire origtmp1605;
	wire origtmp1606;
	wire origtmp1607;
	wire origtmp1608;
	wire origtmp1609;
	wire origtmp1610;
	wire origtmp1611;
	wire origtmp1612;
	wire origtmp1613;
	wire origtmp1614;
	wire origtmp1615;
	wire origtmp1616;
	wire origtmp1617;
	wire origtmp1618;
	wire origtmp1619;
	wire origtmp1620;
	wire origtmp1621;
	wire origtmp1622;
	wire origtmp1623;
	wire origtmp1624;
	wire origtmp1625;
	wire origtmp1626;
	wire origtmp1627;
	wire origtmp1628;
	wire origtmp1629;
	wire origtmp1630;
	wire origtmp1631;
	wire origtmp1632;
	wire origtmp1633;
	wire origtmp1634;
	wire origtmp1635;
	wire origtmp1636;
	wire origtmp1637;
	wire origtmp1638;
	wire origtmp1639;
	wire origtmp1640;
	wire origtmp1641;
	wire origtmp1642;
	wire origtmp1643;
	wire origtmp1644;
	wire origtmp1645;
	wire origtmp1646;
	wire origtmp1647;
	wire origtmp1648;
	wire origtmp1649;
	wire origtmp1650;
	wire origtmp1651;
	wire origtmp1652;
	wire origtmp1653;
	wire origtmp1654;
	wire origtmp1655;
	wire origtmp1656;
	wire origtmp1657;
	wire origtmp1658;
	wire origtmp1659;
	wire origtmp1660;
	wire origtmp1661;
	wire origtmp1662;
	wire origtmp1663;
	wire origtmp1664;
	wire origtmp1665;
	wire origtmp1666;
	wire origtmp1667;
	wire origtmp1668;
	wire origtmp1669;
	wire origtmp1670;
	wire origtmp1671;
	wire origtmp1672;
	wire origtmp1673;
	wire origtmp1674;
	wire origtmp1675;
	wire origtmp1676;
	wire origtmp1677;
	wire origtmp1678;
	wire origtmp1679;
	wire origtmp1680;
	wire origtmp1681;
	wire origtmp1682;
	wire origtmp1683;
	wire origtmp1684;
	wire origtmp1685;
	wire origtmp1686;
	wire origtmp1687;
	wire origtmp1688;
	wire origtmp1689;
	wire origtmp1690;
	wire origtmp1691;
	wire origtmp1692;
	wire origtmp1693;
	wire origtmp1694;
	wire origtmp1695;
	wire origtmp1696;
	wire origtmp1697;
	wire origtmp1698;
	wire origtmp1699;
	wire origtmp1700;
	wire origtmp1701;
	wire origtmp1702;
	wire origtmp1703;
	wire origtmp1704;
	wire origtmp1705;
	wire origtmp1706;
	wire origtmp1707;
	wire origtmp1708;
	wire origtmp1709;
	wire origtmp1710;
	wire origtmp1711;
	wire origtmp1712;
	wire origtmp1713;
	wire origtmp1714;
	wire origtmp1715;
	wire origtmp1716;
	wire origtmp1717;
	wire origtmp1718;
	wire origtmp1719;
	wire origtmp1720;
	wire origtmp1721;
	wire origtmp1722;
	wire origtmp1723;
	wire origtmp1724;
	wire origtmp1725;
	wire origtmp1726;
	wire origtmp1727;
	wire origtmp1728;
	wire origtmp1729;
	wire origtmp1730;
	wire origtmp1731;
	wire origtmp1732;
	wire origtmp1733;
	wire origtmp1734;
	wire origtmp1735;
	wire origtmp1736;
	wire origtmp1737;
	wire origtmp1738;
	wire origtmp1739;
	wire origtmp1740;
	wire origtmp1741;
	wire origtmp1742;
	wire origtmp1743;
	wire origtmp1744;
	wire origtmp1745;
	wire origtmp1746;
	wire origtmp1747;
	wire origtmp1748;
	wire origtmp1749;
	wire origtmp1750;
	wire origtmp1751;
	wire origtmp1752;
	wire origtmp1753;
	wire origtmp1754;
	wire origtmp1755;
	wire origtmp1756;
	wire origtmp1757;
	wire origtmp1758;
	wire origtmp1759;
	wire origtmp1760;
	wire origtmp1761;
	wire origtmp1762;
	wire origtmp1763;
	wire origtmp1764;
	wire origtmp1765;
	wire origtmp1766;
	wire origtmp1767;
	wire origtmp1768;
	wire origtmp1769;
	wire origtmp1770;
	wire origtmp1771;
	wire origtmp1772;
	wire origtmp1773;
	wire origtmp1774;
	wire origtmp1775;
	wire origtmp1776;
	wire origtmp1777;
	wire origtmp1778;
	wire origtmp1779;
	wire origtmp1780;
	wire origtmp1781;
	wire origtmp1782;
	wire origtmp1783;
	wire origtmp1784;
	wire origtmp1785;
	wire origtmp1786;
	wire origtmp1787;
	wire origtmp1788;
	wire origtmp1789;
	wire origtmp1790;
	wire origtmp1791;
	wire origtmp1792;
	wire origtmp1793;
	wire origtmp1794;
	wire origtmp1795;
	wire origtmp1796;
	wire origtmp1797;
	wire origtmp1798;
	wire origtmp1799;
	wire origtmp1800;
	wire origtmp1801;
	wire origtmp1802;
	wire origtmp1803;
	wire origtmp1804;
	wire origtmp1805;
	wire origtmp1806;
	wire origtmp1807;
	wire origtmp1808;
	wire origtmp1809;
	wire origtmp1810;
	wire origtmp1811;
	wire origtmp1812;
	wire origtmp1813;
	wire origtmp1814;
	wire origtmp1815;
	wire origtmp1816;
	wire origtmp1817;
	wire origtmp1818;
	wire origtmp1819;
	wire origtmp1820;
	wire origtmp1821;
	wire origtmp1822;
	wire origtmp1823;
	wire origtmp1824;
	wire origtmp1825;
	wire origtmp1826;
	wire origtmp1827;
	wire origtmp1828;
	wire origtmp1829;
	wire origtmp1830;
	wire origtmp1831;
	wire origtmp1832;
	wire origtmp1833;
	wire origtmp1834;
	wire origtmp1835;
	wire origtmp1836;
	wire origtmp1837;
	wire origtmp1838;
	wire origtmp1839;
	wire origtmp1840;
	wire origtmp1841;
	wire origtmp1842;
	wire origtmp1843;
	wire origtmp1844;
	wire origtmp1845;
	wire origtmp1846;
	wire origtmp1847;
	wire origtmp1848;
	wire origtmp1849;
	wire origtmp1850;
	wire origtmp1851;
	wire origtmp1852;
	wire origtmp1853;
	wire origtmp1854;
	wire origtmp1855;
	wire origtmp1856;
	wire origtmp1857;
	wire origtmp1858;
	wire origtmp1859;
	wire origtmp1860;
	wire origtmp1861;
	wire origtmp1862;
	wire origtmp1863;
	wire origtmp1864;
	wire origtmp1865;
	wire origtmp1866;
	wire origtmp1867;
	wire origtmp1868;
	wire origtmp1869;
	wire origtmp1870;
	wire origtmp1871;
	wire origtmp1872;
	wire origtmp1873;
	wire origtmp1874;
	wire origtmp1875;
	wire origtmp1876;
	wire origtmp1877;
	wire origtmp1878;
	wire origtmp1879;
	wire origtmp1880;
	wire origtmp1881;
	wire origtmp1882;
	wire origtmp1883;
	wire origtmp1884;
	wire origtmp1885;
	wire origtmp1886;
	wire origtmp1887;
	wire origtmp1888;
	wire origtmp1889;
	wire origtmp1890;
	wire origtmp1891;
	wire origtmp1892;
	wire origtmp1893;
	wire origtmp1894;
	wire origtmp1895;
	wire origtmp1896;
	wire origtmp1897;
	wire origtmp1898;
	wire origtmp1899;
	wire origtmp1900;
	wire origtmp1901;
	wire origtmp1902;
	wire origtmp1903;
	wire origtmp1904;
	wire origtmp1905;
	wire origtmp1906;
	wire origtmp1907;
	wire origtmp1908;
	wire origtmp1909;
	wire origtmp1910;
	wire origtmp1911;
	wire origtmp1912;
	wire origtmp1913;
	wire origtmp1914;
	wire origtmp1915;
	wire origtmp1916;
	wire origtmp1917;
	wire origtmp1918;
	wire origtmp1919;
	wire origtmp1920;
	wire origtmp1921;
	wire origtmp1922;
	wire origtmp1923;
	wire origtmp1924;
	wire origtmp1925;
	wire origtmp1926;
	wire origtmp1927;
	wire origtmp1928;
	wire origtmp1929;
	wire origtmp1930;
	wire origtmp1931;
	wire origtmp1932;
	wire origtmp1933;
	wire origtmp1934;
	wire origtmp1935;
	wire origtmp1936;
	wire origtmp1937;
	wire origtmp1938;
	wire origtmp1939;
	wire origtmp1940;
	wire origtmp1941;
	wire origtmp1942;
	wire origtmp1943;
	wire origtmp1944;
	wire origtmp1945;
	wire origtmp1946;
	wire origtmp1947;
	wire origtmp1948;
	wire origtmp1949;
	wire origtmp1950;
	wire origtmp1951;
	wire origtmp1952;
	wire origtmp1953;
	wire origtmp1954;
	wire origtmp1955;
	wire origtmp1956;
	wire origtmp1957;
	wire origtmp1958;
	wire origtmp1959;
	wire origtmp1960;
	wire origtmp1961;
	wire origtmp1962;
	wire origtmp1963;
	wire origtmp1964;
	wire origtmp1965;
	wire origtmp1966;
	wire origtmp1967;
	wire origtmp1968;
	wire origtmp1969;
	wire origtmp1970;
	wire origtmp1971;
	wire origtmp1972;
	wire origtmp1973;
	wire origtmp1974;
	wire origtmp1975;
	wire origtmp1976;
	wire origtmp1977;
	wire origtmp1978;
	wire origtmp1979;
	wire origtmp1980;
	wire origtmp1981;
	wire origtmp1982;
	wire origtmp1983;
	wire origtmp1984;
	wire origtmp1985;
	wire origtmp1986;
	wire origtmp1987;
	wire origtmp1988;
	wire origtmp1989;
	wire origtmp1990;
	wire origtmp1991;
	wire origtmp1992;
	wire origtmp1993;
	wire origtmp1994;
	wire origtmp1995;
	wire origtmp1996;
	wire origtmp1997;
	wire origtmp1998;
	wire origtmp1999;
	wire origtmp2000;
	wire origtmp2001;
	wire origtmp2002;
	wire origtmp2003;
	wire origtmp2004;
	wire origtmp2005;
	wire origtmp2006;
	wire origtmp2007;
	wire origtmp2008;
	wire origtmp2009;
	wire origtmp2010;
	wire origtmp2011;
	wire origtmp2012;
	wire origtmp2013;
	wire origtmp2014;
	wire origtmp2015;
	wire origtmp2016;
	wire origtmp2017;
	wire origtmp2018;
	wire origtmp2019;
	wire origtmp2020;
	wire origtmp2021;
	wire origtmp2022;
	wire origtmp2023;
	wire origtmp2024;
	wire origtmp2025;
	wire origtmp2026;
	wire origtmp2027;
	wire origtmp2028;
	wire origtmp2029;
	wire origtmp2030;
	wire origtmp2031;
	wire origtmp2032;
	wire origtmp2033;
	wire origtmp2034;
	wire origtmp2035;
	wire origtmp2036;
	wire origtmp2037;
	wire origtmp2038;
	wire origtmp2039;
	wire origtmp2040;
	wire origtmp2041;
	wire origtmp2042;
	wire origtmp2043;
	wire origtmp2044;
	wire origtmp2045;
	wire origtmp2046;
	wire origtmp2047;
	wire origtmp2048;
	wire origtmp2049;
	wire origtmp2050;
	wire origtmp2051;
	wire origtmp2052;
	wire origtmp2053;
	wire origtmp2054;
	wire origtmp2055;
	wire origtmp2056;
	wire origtmp2057;
	wire origtmp2058;
	wire origtmp2059;
	wire origtmp2060;
	wire origtmp2061;
	wire origtmp2062;
	wire origtmp2063;
	wire origtmp2064;
	wire origtmp2065;
	wire origtmp2066;
	wire origtmp2067;
	wire origtmp2068;
	wire origtmp2069;
	wire origtmp2070;
	wire origtmp2071;
	wire origtmp2072;
	wire origtmp2073;
	wire origtmp2074;
	wire origtmp2075;
	wire origtmp2076;
	wire origtmp2077;
	wire origtmp2078;
	wire origtmp2079;
	wire origtmp2080;
	wire origtmp2081;
	wire origtmp2082;
	wire origtmp2083;
	wire origtmp2084;
	wire origtmp2085;
	wire origtmp2086;
	wire origtmp2087;
	wire origtmp2088;
	wire origtmp2089;
	wire origtmp2090;
	wire origtmp2091;
	wire origtmp2092;
	wire origtmp2093;
	wire origtmp2094;
	wire origtmp2095;
	wire origtmp2096;
	wire origtmp2097;
	wire origtmp2098;
	wire origtmp2099;
	wire origtmp2100;
	wire origtmp2101;
	wire origtmp2102;
	wire origtmp2103;
	wire origtmp2104;
	wire origtmp2105;
	wire origtmp2106;
	wire origtmp2107;
	wire origtmp2108;
	wire origtmp2109;
	wire origtmp2110;
	wire origtmp2111;
	wire origtmp2112;
	wire origtmp2113;
	wire origtmp2114;
	wire origtmp2115;
	wire origtmp2116;
	wire origtmp2117;
	wire origtmp2118;
	wire origtmp2119;
	wire origtmp2120;
	wire origtmp2121;
	wire origtmp2122;
	wire origtmp2123;
	wire origtmp2124;
	wire origtmp2125;
	wire origtmp2126;
	wire origtmp2127;
	wire origtmp2128;
	wire origtmp2129;
	wire origtmp2130;
	wire origtmp2131;
	wire origtmp2132;
	wire origtmp2133;
	wire origtmp2134;
	wire origtmp2135;
	wire origtmp2136;
	wire origtmp2137;
	wire origtmp2138;
	wire origtmp2139;
	wire origtmp2140;
	wire origtmp2141;
	wire origtmp2142;
	wire origtmp2143;
	wire origtmp2144;
	wire origtmp2145;
	wire origtmp2146;
	wire origtmp2147;
	wire origtmp2148;
	wire origtmp2149;
	wire origtmp2150;
	wire origtmp2151;
	wire origtmp2152;
	wire origtmp2153;
	wire origtmp2154;
	wire origtmp2155;
	wire origtmp2156;
	wire origtmp2157;
	wire origtmp2158;
	wire origtmp2159;
	wire origtmp2160;
	wire origtmp2161;
	wire origtmp2162;
	wire origtmp2163;
	wire origtmp2164;
	wire origtmp2165;
	wire origtmp2166;
	wire origtmp2167;
	wire origtmp2168;
	wire origtmp2169;
	wire origtmp2170;
	wire origtmp2171;
	wire origtmp2172;
	wire origtmp2173;
	wire origtmp2174;
	wire origtmp2175;
	wire origtmp2176;
	wire origtmp2177;
	wire origtmp2178;
	wire origtmp2179;
	wire origtmp2180;
	wire origtmp2181;
	wire origtmp2182;
	wire origtmp2183;
	wire origtmp2184;
	wire origtmp2185;
	wire origtmp2186;
	wire origtmp2187;
	wire origtmp2188;
	wire origtmp2189;
	wire origtmp2190;
	wire origtmp2191;
	wire origtmp2192;
	wire origtmp2193;
	wire origtmp2194;
	wire origtmp2195;
	wire origtmp2196;
	wire origtmp2197;
	wire origtmp2198;
	wire origtmp2199;
	wire origtmp2200;
	wire origtmp2201;
	wire origtmp2202;
	wire origtmp2203;
	wire origtmp2204;
	wire origtmp2205;
	wire origtmp2206;
	wire origtmp2207;
	wire origtmp2208;
	wire origtmp2209;
	wire origtmp2210;
	wire origtmp2211;
	wire origtmp2212;
	wire origtmp2213;
	wire origtmp2214;
	wire origtmp2215;
	wire origtmp2216;
	wire origtmp2217;
	wire origtmp2218;
	wire origtmp2219;
	wire origtmp2220;
	wire origtmp2221;
	wire origtmp2222;
	wire origtmp2223;
	wire origtmp2224;
	wire origtmp2225;
	wire origtmp2226;
	wire origtmp2227;
	wire origtmp2228;
	wire origtmp2229;
	wire origtmp2230;
	wire origtmp2231;
	wire origtmp2232;
	wire origtmp2233;
	wire origtmp2234;
	wire origtmp2235;
	wire origtmp2236;
	wire origtmp2237;
	wire origtmp2238;
	wire origtmp2239;
	wire origtmp2240;
	wire origtmp2241;
	wire origtmp2242;
	wire origtmp2243;
	wire origtmp2244;
	wire origtmp2245;
	wire origtmp2246;
	wire origtmp2247;
	wire origtmp2248;
	wire origtmp2249;
	wire origtmp2250;
	wire origtmp2251;
	wire origtmp2252;
	wire origtmp2253;
	wire origtmp2254;
	wire origtmp2255;
	wire origtmp2256;
	assign out[92] = origtmp228 & origtmp229;
	assign out[134] = origtmp331 | 1'b1;
	assign origtmp2032 = in[1365] | in[994];
	assign out[219] = origtmp546;
	assign origtmp966 = origtmp967 & origtmp965;
	assign origtmp1472 = origtmp1373 | origtmp1722;
	assign origtmp1015 = in[24] ^ in[24];
	assign origtmp36 = in[749] & origtmp35;
	assign origtmp1976 = origtmp1895 ^ in[1071];
	assign origtmp1048 = origtmp1049 | origtmp1050;
	assign out[278] = origtmp699 | origtmp700;
	assign out[64] = origtmp162 & origtmp160;
	assign origtmp2154 = origtmp2080 & in[1279];
	assign origtmp725 = origtmp724 ^ in[220];
	assign out[80] = 1'b1 | 1'b0;
	assign out[300] = origtmp753;
	assign origtmp408 = 1'b0 | 1'b1;
	assign origtmp1074 = in[1309] & 1'b0;
	assign origtmp401 = origtmp398 ^ origtmp402;
	assign out[165] = origtmp413 ^ in[1302];
	assign origtmp2017 = in[671] & in[155];
	assign origtmp1557 = origtmp1638 & origtmp1267;
	assign origtmp1690 = in[1163] | origtmp1260;
	assign out[466] = origtmp1168 | origtmp1168;
	assign origtmp1881 = origtmp2029 & in[125];
	assign origtmp617 = in[131] | 1'b0;
	assign out[461] = origtmp1156 ^ in[252];
	assign origtmp2232 = in[473] & in[714];
	assign origtmp1602 = in[518] | in[1042];
	assign origtmp762 = origtmp763 ^ in[695];
	assign out[148] = origtmp366 ^ in[1107];
	assign origtmp1192 = in[332] & 1'b0;
	assign origtmp2182 = origtmp2122 ^ origtmp1247;
	assign out[206] = in[1394];
	assign origtmp615 = in[258] | in[650];
	assign origtmp1487 = in[1154] & origtmp2191;
	assign origtmp474 = ~1'b0;
	assign origtmp53 = ~in[1101];
	assign origtmp1960 = origtmp1950 ^ origtmp1969;
	assign out[170] = origtmp425 | origtmp425;
	assign origtmp949 = origtmp950 & origtmp950;
	assign origtmp390 = origtmp388 & in[9];
	assign origtmp2231 = in[873] & origtmp1528;
	assign out[222] = origtmp556 & 1'b0;
	assign origtmp2101 = in[995] | in[1450];
	assign origtmp1091 = 1'b0 & 1'b1;
	assign out[336] = origtmp839 & 1'b0;
	assign origtmp1255 = in[1280] | in[902];
	assign origtmp1157 = ~1'b1;
	assign origtmp1240 = origtmp1237 ^ 1'b0;
	assign origtmp838 = in[986];
	assign origtmp485 = 1'b1 & 1'b0;
	assign origtmp740 = in[809] & in[799];
	assign origtmp606 = 1'b0 | origtmp605;
	assign origtmp356 = 1'b0 & origtmp358;
	assign origtmp858 = origtmp857 ^ in[425];
	assign origtmp1761 = origtmp2019 & origtmp1955;
	assign origtmp172 = 1'b0;
	assign origtmp591 = origtmp592 | 1'b0;
	assign origtmp773 = 1'b0 ^ origtmp772;
	assign out[267] = origtmp666 ^ origtmp667;
	assign out[205] = ~1'b1;
	assign origtmp1998 = in[1248] & in[303];
	assign origtmp1644 = origtmp1873 ^ origtmp1288;
	assign origtmp2081 = origtmp1912 | origtmp1750;
	assign out[121] = origtmp300 | in[1402];
	assign out[493] = 1'b0 | origtmp1232;
	assign origtmp492 = origtmp494 | 1'b1;
	assign origtmp760 = ~1'b0;
	assign origtmp1997 = in[1373] ^ in[1220];
	assign out[228] = origtmp573 | origtmp574;
	assign out[99] = 1'b0 | origtmp249;
	assign origtmp1700 = origtmp1591 ^ origtmp1268;
	assign origtmp1981 = in[1086] & in[1214];
	assign origtmp1465 = origtmp1585 ^ origtmp1664;
	assign origtmp620 = origtmp621 & in[1005];
	assign out[286] = ~origtmp725;
	assign origtmp931 = in[33] & 1'b0;
	assign origtmp1616 = in[778] ^ origtmp2014;
	assign out[137] = origtmp337 | origtmp336;
	assign origtmp859 = 1'b1;
	assign origtmp291 = 1'b1 ^ origtmp289;
	assign origtmp1001 = 1'b1 ^ 1'b0;
	assign origtmp1092 = in[1361] & origtmp1095;
	assign out[428] = 1'b0 | origtmp1064;
	assign out[287] = origtmp727 & origtmp726;
	assign origtmp524 = 1'b1 | origtmp522;
	assign origtmp1350 = origtmp1856 ^ in[397];
	assign origtmp548 = 1'b0;
	assign origtmp718 = origtmp720 ^ origtmp719;
	assign origtmp876 = origtmp874 | origtmp874;
	assign origtmp588 = ~1'b0;
	assign origtmp815 = ~1'b1;
	assign out[7] = in[1474] & origtmp11;
	assign origtmp1825 = origtmp1545 ^ in[992];
	assign out[88] = origtmp221 & 1'b1;
	assign origtmp711 = 1'b1 ^ in[697];
	assign out[478] = origtmp1201 & origtmp1202;
	assign origtmp1332 = origtmp1729 ^ origtmp1872;
	assign origtmp1794 = in[1261] ^ in[45];
	assign origtmp386 = ~origtmp390;
	assign origtmp361 = 1'b1 & in[1143];
	assign origtmp2131 = in[769] & origtmp1627;
	assign origtmp1412 = in[381] ^ in[581];
	assign origtmp1680 = in[1203] ^ in[242];
	assign origtmp11 = origtmp10;
	assign origtmp349 = in[630] ^ origtmp350;
	assign origtmp2121 = in[700] ^ in[1176];
	assign origtmp272 = in[1089] ^ in[1089];
	assign origtmp2166 = in[46] & in[333];
	assign origtmp1326 = in[698] ^ origtmp1926;
	assign origtmp748 = origtmp747 | in[285];
	assign origtmp1460 = in[363] | in[840];
	assign out[299] = origtmp749 & origtmp748;
	assign origtmp288 = in[511] | origtmp290;
	assign origtmp1438 = origtmp1776 | origtmp1654;
	assign out[345] = origtmp858;
	assign out[366] = in[1134] & origtmp905;
	assign origtmp1349 = in[707] ^ origtmp1700;
	assign origtmp358 = in[390] ^ 1'b0;
	assign origtmp1481 = in[465] ^ origtmp1784;
	assign origtmp210 = 1'b0 & origtmp211;
	assign origtmp1210 = in[649] ^ in[1400];
	assign out[33] = origtmp87 ^ origtmp86;
	assign origtmp157 = ~in[516];
	assign origtmp1466 = origtmp1595 ^ origtmp1931;
	assign origtmp340 = in[1335];
	assign out[460] = 1'b0;
	assign origtmp1060 = origtmp1061 & 1'b0;
	assign origtmp1966 = origtmp1774 | origtmp1691;
	assign origtmp793 = in[1234] & 1'b0;
	assign origtmp1941 = origtmp1506 ^ in[1155];
	assign origtmp1936 = origtmp1878 ^ origtmp1303;
	assign origtmp1410 = origtmp1248 ^ origtmp2103;
	assign origtmp339 = in[1335] & 1'b1;
	assign out[168] = origtmp414 | origtmp416;
	assign origtmp241 = origtmp238 | in[1293];
	assign origtmp1257 = origtmp2013 | origtmp1975;
	assign origtmp461 = in[715] | origtmp459;
	assign out[220] = origtmp550 & in[488];
	assign origtmp566 = in[1142] ^ 1'b1;
	assign origtmp396 = in[1167] & 1'b1;
	assign origtmp509 = in[922];
	assign origtmp2142 = origtmp1834 | in[1063];
	assign out[86] = origtmp215 | origtmp212;
	assign origtmp1140 = 1'b0;
	assign origtmp1377 = origtmp1599 & origtmp1287;
	assign origtmp1718 = in[1024] | origtmp1484;
	assign origtmp2132 = origtmp1544 & origtmp1606;
	assign origtmp975 = 1'b0 & 1'b1;
	assign origtmp1411 = origtmp1705 | origtmp1546;
	assign origtmp2227 = origtmp1504 | origtmp1709;
	assign origtmp1314 = in[43] ^ origtmp1847;
	assign origtmp1898 = in[746] ^ in[1325];
	assign origtmp2164 = origtmp2176 & origtmp1265;
	assign origtmp959 = 1'b1 & in[590];
	assign origtmp2183 = in[1087] & in[621];
	assign origtmp1067 = 1'b0 ^ origtmp1066;
	assign origtmp1233 = in[754] | in[627];
	assign origtmp2004 = in[886] & in[280];
	assign origtmp1391 = origtmp1538 & origtmp1986;
	assign out[140] = origtmp346 & in[1044];
	assign origtmp1322 = in[535] ^ in[344];
	assign out[322] = origtmp801 & origtmp799;
	assign origtmp1590 = in[358] ^ in[1313];
	assign origtmp121 = 1'b0 | in[83];
	assign origtmp912 = 1'b1 | 1'b1;
	assign origtmp985 = ~1'b1;
	assign out[254] = origtmp632 | origtmp632;
	assign origtmp2241 = in[507] ^ origtmp1849;
	assign origtmp1143 = origtmp1145 & in[328];
	assign origtmp501 = 1'b0 ^ 1'b1;
	assign origtmp467 = in[1269] | origtmp468;
	assign out[203] = in[800] ^ 1'b1;
	assign origtmp334 = origtmp333;
	assign origtmp495 = origtmp496 & origtmp496;
	assign out[273] = 1'b0 | origtmp683;
	assign origtmp235 = origtmp236 | in[1357];
	assign origtmp369 = in[1387] | 1'b1;
	assign out[174] = origtmp439 ^ origtmp437;
	assign origtmp1030 = 1'b1;
	assign origtmp733 = ~1'b0;
	assign out[214] = origtmp530 | origtmp528;
	assign origtmp1373 = origtmp2085 ^ in[1205];
	assign origtmp545 = 1'b0 & 1'b0;
	assign origtmp1246 = origtmp1410 | in[903];
	assign origtmp1884 = origtmp2231 | in[834];
	assign out[435] = in[896] & 1'b1;
	assign origtmp1375 = origtmp1925 ^ origtmp1636;
	assign origtmp1371 = in[1121] | origtmp1311;
	assign origtmp687 = 1'b0;
	assign origtmp676 = in[202] | 1'b1;
	assign origtmp1812 = in[113] ^ in[958];
	assign origtmp243 = origtmp242 | origtmp245;
	assign origtmp819 = in[210] | 1'b1;
	assign origtmp698 = origtmp697 | in[976];
	assign origtmp1561 = origtmp2048 | origtmp1633;
	assign origtmp1445 = origtmp1598 | origtmp1294;
	assign origtmp1254 = origtmp1976 ^ origtmp1646;
	assign origtmp643 = origtmp640 | in[7];
	assign origtmp1301 = origtmp2186 ^ origtmp1893;
	assign origtmp1840 = in[311] | origtmp1344;
	assign origtmp47 = origtmp45 ^ origtmp43;
	assign out[439] = in[1178] & origtmp1086;
	assign origtmp44 = origtmp47 & origtmp46;
	assign out[253] = in[380] | origtmp631;
	assign origtmp1977 = origtmp1626 & in[406];
	assign origtmp1292 = origtmp1823 | in[965];
	assign origtmp1390 = origtmp2004 | in[1446];
	assign out[337] = origtmp840 & 1'b0;
	assign origtmp1129 = origtmp1127;
	assign origtmp1151 = origtmp1153 & 1'b0;
	assign origtmp1462 = in[246] & origtmp1372;
	assign out[146] = origtmp360 & origtmp361;
	assign origtmp1736 = origtmp2183 | in[779];
	assign origtmp1576 = origtmp2167 | in[836];
	assign origtmp1532 = origtmp1286 & in[951];
	assign origtmp1702 = origtmp1884 ^ in[1105];
	assign origtmp1334 = origtmp1537 | origtmp1262;
	assign origtmp1333 = in[1009] & in[1128];
	assign origtmp1594 = in[1281] ^ in[224];
	assign origtmp2185 = origtmp1594 | in[114];
	assign origtmp1845 = in[1316] & origtmp1831;
	assign out[356] = origtmp889 & origtmp889;
	assign origtmp1093 = 1'b0 | 1'b0;
	assign origtmp1339 = in[1452] & origtmp1394;
	assign origtmp95 = 1'b0;
	assign origtmp1426 = in[121] | in[1125];
	assign out[25] = origtmp67 | origtmp65;
	assign origtmp1567 = origtmp2092 | in[472];
	assign origtmp2172 = in[1223] & in[1120];
	assign out[341] = origtmp851 & origtmp850;
	assign origtmp2107 = origtmp1837 | origtmp1686;
	assign origtmp38 = 1'b0 & origtmp37;
	assign origtmp1771 = origtmp1892 & in[694];
	assign origtmp597 = in[1236] ^ origtmp595;
	assign origtmp1531 = in[1443] ^ origtmp1608;
	assign origtmp772 = 1'b0;
	assign origtmp267 = 1'b1 | origtmp266;
	assign origtmp752 = ~origtmp754;
	assign origtmp1753 = in[913] | in[237];
	assign origtmp1580 = in[61] & in[688];
	assign origtmp1883 = in[1053] & in[1160];
	assign origtmp403 = origtmp404 ^ 1'b0;
	assign out[331] = ~origtmp825;
	assign origtmp465 = in[681] & origtmp464;
	assign origtmp268 = 1'b1 ^ origtmp269;
	assign origtmp1253 = in[312] | in[1252];
	assign origtmp791 = origtmp790 | origtmp790;
	assign origtmp729 = origtmp730;
	assign origtmp204 = 1'b1 & origtmp203;
	assign origtmp1502 = in[92] & origtmp1778;
	assign origtmp944 = origtmp946 ^ in[1350];
	assign out[418] = 1'b1 | origtmp1030;
	assign origtmp2011 = origtmp1357 | origtmp1775;
	assign origtmp1066 = 1'b0;
	assign out[473] = origtmp1189 ^ origtmp1191;
	assign origtmp837 = origtmp838 ^ 1'b0;
	assign origtmp1957 = origtmp2060 | origtmp1423;
	assign origtmp1823 = origtmp1930 ^ origtmp1885;
	assign out[450] = origtmp1120 & origtmp1123;
	assign origtmp662 = origtmp665 | origtmp663;
	assign origtmp738 = in[500];
	assign origtmp1926 = in[1410] ^ in[1068];
	assign origtmp97 = ~1'b0;
	assign out[32] = origtmp82 | origtmp84;
	assign origtmp2076 = in[830] | origtmp1602;
	assign origtmp164 = 1'b0 | in[403];
	assign out[455] = origtmp1138 ^ origtmp1141;
	assign origtmp127 = 1'b0 ^ 1'b0;
	assign out[302] = origtmp759 | origtmp759;
	assign origtmp834 = origtmp835 | 1'b0;
	assign out[386] = origtmp955 | origtmp953;
	assign out[495] = in[159] | 1'b1;
	assign origtmp2256 = origtmp1558 | origtmp2251;
	assign origtmp1814 = in[943] | origtmp1735;
	assign out[320] = origtmp795 ^ 1'b1;
	assign out[127] = in[1268] ^ origtmp320;
	assign origtmp775 = in[810] & in[1179];
	assign origtmp1228 = in[79] & origtmp1226;
	assign origtmp2116 = in[404] ^ in[1130];
	assign origtmp214 = ~origtmp213;
	assign out[275] = origtmp691 & origtmp690;
	assign origtmp737 = ~in[500];
	assign origtmp365 = 1'b1 & origtmp362;
	assign origtmp1492 = origtmp1897 & origtmp1906;
	assign out[268] = origtmp668 ^ origtmp668;
	assign origtmp1296 = in[1151] ^ origtmp2234;
	assign origtmp2028 = in[531] | origtmp1413;
	assign origtmp2043 = origtmp1397 ^ in[1409];
	assign out[5] = 1'b0;
	assign out[84] = origtmp207 | origtmp207;
	assign origtmp1446 = in[31] | origtmp1507;
	assign origtmp336 = origtmp340 ^ origtmp338;
	assign origtmp1018 = 1'b0 ^ origtmp1017;
	assign out[391] = 1'b1 | origtmp966;
	assign origtmp145 = origtmp144 | origtmp146;
	assign origtmp1779 = in[227] ^ in[1419];
	assign origtmp1286 = in[1441] | in[577];
	assign origtmp458 = origtmp455 | origtmp456;
	assign out[139] = in[221] ^ origtmp342;
	assign origtmp2159 = in[1000] ^ origtmp2245;
	assign origtmp1423 = in[996] ^ in[596];
	assign origtmp1583 = origtmp2215 ^ in[352];
	assign out[262] = 1'b1 ^ in[593];
	assign origtmp1278 = in[1140] & origtmp1953;
	assign origtmp1604 = origtmp1568 ^ in[1287];
	assign origtmp479 = origtmp478;
	assign origtmp2151 = in[1290] | origtmp1688;
	assign out[113] = origtmp286 & 1'b1;
	assign origtmp277 = in[387] | origtmp276;
	assign origtmp1660 = origtmp1734 ^ in[1091];
	assign origtmp982 = origtmp986 & 1'b1;
	assign origtmp1648 = origtmp1909 | origtmp1850;
	assign origtmp1470 = in[863] & in[134];
	assign origtmp1242 = in[1385] ^ in[65];
	assign origtmp1499 = in[88] | in[1482];
	assign origtmp1008 = ~in[802];
	assign out[459] = origtmp1154 | origtmp1151;
	assign origtmp1552 = in[683] & in[732];
	assign origtmp2175 = origtmp1252 ^ in[1035];
	assign origtmp1944 = in[268] ^ origtmp1604;
	assign origtmp941 = ~in[347];
	assign origtmp1638 = in[878] ^ in[782];
	assign origtmp1928 = in[1030] ^ in[1270];
	assign out[289] = origtmp732 & origtmp734;
	assign origtmp1176 = 1'b1 | in[971];
	assign out[242] = ~origtmp603;
	assign origtmp678 = origtmp682 ^ origtmp681;
	assign origtmp134 = origtmp136 | origtmp132;
	assign origtmp101 = origtmp100 & origtmp100;
	assign out[39] = origtmp102 ^ 1'b0;
	assign origtmp3 = ~1'b1;
	assign out[129] = in[1241] & 1'b1;
	assign origtmp742 = 1'b1 | in[809];
	assign origtmp1315 = in[119] | in[1033];
	assign out[469] = in[600] ^ origtmp1177;
	assign origtmp2113 = origtmp1640 ^ in[819];
	assign origtmp450 = ~1'b1;
	assign origtmp2187 = origtmp1692 | in[442];
	assign origtmp2250 = origtmp2242 & origtmp1459;
	assign origtmp1862 = in[314] & in[300];
	assign origtmp1174 = 1'b1 | origtmp1175;
	assign origtmp1497 = in[467] ^ origtmp1520;
	assign origtmp822 = in[936] | origtmp819;
	assign origtmp58 = 1'b0;
	assign out[231] = origtmp580 ^ in[152];
	assign origtmp828 = origtmp830 & in[833];
	assign origtmp604 = origtmp601;
	assign origtmp1634 = origtmp1533 ^ in[954];
	assign origtmp881 = origtmp878 & origtmp878;
	assign origtmp1890 = origtmp2112 & in[1330];
	assign out[412] = origtmp1011 | origtmp1011;
	assign origtmp1324 = origtmp1275 & in[1187];
	assign origtmp1031 = 1'b1 & in[1123];
	assign origtmp1136 = 1'b1 ^ in[1383];
	assign origtmp5 = in[1456] ^ 1'b1;
	assign origtmp572 = origtmp570 ^ origtmp569;
	assign out[380] = origtmp936;
	assign origtmp2045 = origtmp1431 ^ origtmp1861;
	assign origtmp919 = in[194] | in[168];
	assign origtmp1206 = in[1497] ^ 1'b0;
	assign origtmp265 = 1'b0 | 1'b1;
	assign origtmp1504 = in[44] ^ in[376];
	assign origtmp849 = 1'b0 & in[1328];
	assign out[431] = origtmp1070 | origtmp1072;
	assign origtmp1399 = in[71] & in[192];
	assign out[295] = in[947] | 1'b1;
	assign origtmp1542 = in[392] | origtmp1811;
	assign origtmp111 = in[1278] | 1'b1;
	assign origtmp641 = 1'b1 & 1'b0;
	assign origtmp1972 = origtmp1500 | in[1285];
	assign origtmp1584 = origtmp1471 | origtmp1666;
	assign origtmp205 = 1'b0 | origtmp204;
	assign origtmp522 = in[444] & origtmp521;
	assign origtmp1992 = in[181] | origtmp1519;
	assign origtmp570 = 1'b0;
	assign origtmp460 = 1'b1 & origtmp462;
	assign origtmp308 = ~origtmp307;
	assign out[265] = origtmp660 & origtmp659;
	assign origtmp1040 = in[122] & in[1311];
	assign origtmp1194 = in[332] | origtmp1192;
	assign origtmp46 = 1'b0 | 1'b0;
	assign origtmp1819 = origtmp1306 ^ origtmp2182;
	assign origtmp2102 = origtmp1529 | origtmp1745;
	assign origtmp156 = origtmp155 | origtmp153;
	assign origtmp42 = in[1314] & in[1314];
	assign origtmp1916 = origtmp1716 | in[426];
	assign origtmp902 = origtmp904 ^ origtmp904;
	assign origtmp1297 = origtmp2003 | in[609];
	assign origtmp1467 = in[679] & in[625];
	assign out[40] = origtmp104 ^ in[933];
	assign origtmp1946 = in[604] & in[720];
	assign origtmp979 = in[1039];
	assign origtmp686 = 1'b1 | 1'b1;
	assign origtmp1887 = origtmp2180 | origtmp1378;
	assign origtmp456 = 1'b0;
	assign origtmp55 = origtmp58 | origtmp56;
	assign origtmp420 = origtmp421 ^ origtmp421;
	assign out[166] = 1'b1 | 1'b0;
	assign origtmp457 = in[885] | origtmp456;
	assign origtmp1084 = ~origtmp1082;
	assign origtmp999 = 1'b1;
	assign origtmp777 = 1'b1 | in[810];
	assign origtmp1646 = in[934] & origtmp2171;
	assign origtmp1754 = in[236] ^ in[1181];
	assign origtmp436 = in[539] | origtmp432;
	assign origtmp503 = origtmp499 ^ in[549];
	assign origtmp1514 = origtmp1900 & in[1487];
	assign origtmp256 = 1'b0 ^ origtmp254;
	assign origtmp409 = origtmp408 ^ 1'b0;
	assign origtmp1525 = origtmp1694 | origtmp2046;
	assign origtmp304 = origtmp306 & origtmp305;
	assign origtmp1457 = origtmp1282 | origtmp2143;
	assign origtmp1805 = in[164] | in[1036];
	assign out[18] = origtmp44 ^ 1'b0;
	assign origtmp2092 = origtmp1653 | origtmp1419;
	assign origtmp426 = 1'b0 & in[35];
	assign origtmp248 = origtmp250 ^ origtmp250;
	assign origtmp1515 = in[165] & origtmp1478;
	assign origtmp411 = ~in[949];
	assign origtmp2195 = in[1199] ^ in[1245];
	assign origtmp1923 = origtmp2110 & origtmp1810;
	assign origtmp1213 = origtmp1211 | origtmp1210;
	assign origtmp275 = origtmp274 & in[387];
	assign origtmp1238 = origtmp1237;
	assign origtmp1562 = origtmp1813 & in[39];
	assign origtmp198 = origtmp200 | in[963];
	assign origtmp1758 = in[745] ^ in[433];
	assign origtmp1688 = origtmp2244 & in[684];
	assign origtmp137 = ~in[808];
	assign origtmp996 = in[1169] | in[47];
	assign origtmp526 = 1'b1 & 1'b0;
	assign origtmp2082 = origtmp2133 ^ origtmp2134;
	assign origtmp960 = in[1271] ^ in[230];
	assign out[312] = origtmp782 | origtmp781;
	assign out[434] = origtmp1078 & origtmp1080;
	assign origtmp942 = origtmp945 | origtmp944;
	assign origtmp923 = 1'b0 & 1'b0;
	assign origtmp544 = 1'b1 | 1'b0;
	assign origtmp394 = in[583] & in[709];
	assign origtmp1433 = origtmp1822 ^ origtmp1634;
	assign out[378] = origtmp932 & origtmp934;
	assign origtmp674 = origtmp676 | 1'b0;
	assign origtmp805 = 1'b0;
	assign origtmp565 = ~origtmp564;
	assign origtmp1909 = in[723] | in[821];
	assign origtmp1566 = in[1244] & in[1378];
	assign origtmp338 = 1'b0 ^ 1'b0;
	assign origtmp1207 = in[1497];
	assign origtmp1775 = in[850] ^ in[716];
	assign out[15] = origtmp33 & in[749];
	assign origtmp1942 = origtmp1843 | in[1451];
	assign origtmp444 = 1'b0;
	assign origtmp1516 = in[1249] ^ in[631];
	assign out[283] = origtmp714 ^ origtmp717;
	assign out[398] = origtmp987 | in[1413];
	assign origtmp790 = 1'b0 | 1'b0;
	assign origtmp561 = origtmp557;
	assign out[115] = in[1164] | origtmp292;
	assign origtmp1408 = origtmp1281 | origtmp1456;
	assign out[55] = origtmp135 | origtmp134;
	assign origtmp706 = ~origtmp705;
	assign origtmp534 = in[1415] | 1'b0;
	assign origtmp1752 = origtmp1309 & origtmp1904;
	assign origtmp1204 = in[1298] ^ 1'b1;
	assign origtmp2236 = in[665] & origtmp1874;
	assign out[117] = 1'b1 & 1'b0;
	assign out[468] = origtmp1174 | in[971];
	assign origtmp976 = ~origtmp974;
	assign origtmp962 = origtmp961;
	assign origtmp2083 = in[1078] | in[1388];
	assign origtmp2190 = origtmp1659 | origtmp1455;
	assign origtmp2243 = in[37] | in[1431];
	assign origtmp45 = 1'b0 & in[930];
	assign origtmp1767 = in[32] & in[550];
	assign origtmp1344 = in[393] | origtmp1914;
	assign out[224] = ~origtmp565;
	assign origtmp452 = in[185] & in[185];
	assign origtmp2128 = origtmp1690 ^ origtmp1327;
	assign origtmp523 = origtmp524 | origtmp522;
	assign origtmp537 = origtmp540 | 1'b0;
	assign origtmp2219 = origtmp1552 ^ origtmp2097;
	assign origtmp564 = in[1142] & origtmp562;
	assign out[479] = 1'b1;
	assign origtmp223 = 1'b0 ^ origtmp224;
	assign origtmp89 = 1'b1;
	assign origtmp973 = origtmp975 & origtmp975;
	assign origtmp897 = origtmp899 | origtmp899;
	assign origtmp1945 = origtmp1656 | origtmp1481;
	assign origtmp1202 = ~origtmp1200;
	assign origtmp68 = in[952];
	assign origtmp1239 = origtmp1240 & in[474];
	assign origtmp1216 = origtmp1217 & 1'b0;
	assign origtmp1661 = in[1353] | in[1404];
	assign origtmp464 = in[842] | 1'b1;
	assign origtmp1451 = in[245] & in[1006];
	assign origtmp1319 = origtmp2214 ^ origtmp1447;
	assign origtmp120 = origtmp122 & 1'b0;
	assign origtmp647 = 1'b0 | 1'b1;
	assign out[482] = origtmp1209 | origtmp1209;
	assign origtmp2053 = origtmp2091 ^ in[939];
	assign out[135] = origtmp332;
	assign origtmp610 = 1'b0 & in[57];
	assign origtmp1831 = in[794] & in[357];
	assign origtmp704 = 1'b1;
	assign origtmp991 = origtmp993 ^ in[1020];
	assign origtmp2072 = in[887] & origtmp2030;
	assign origtmp953 = ~1'b0;
	assign origtmp1694 = origtmp1668 & origtmp2095;
	assign origtmp1697 = origtmp1689 & in[508];
	assign origtmp1494 = in[335] & in[494];
	assign origtmp2069 = in[1491] ^ in[1082];
	assign out[46] = 1'b1 ^ 1'b0;
	assign origtmp2224 = origtmp2150 ^ origtmp1246;
	assign origtmp868 = origtmp870 | origtmp870;
	assign origtmp1523 = origtmp1428 & in[696];
	assign origtmp1854 = origtmp1902 ^ origtmp2096;
	assign origtmp847 = 1'b0 | 1'b1;
	assign origtmp366 = in[1107] | in[1107];
	assign origtmp1991 = origtmp1657 & origtmp1848;
	assign origtmp629 = origtmp627 ^ in[1460];
	assign origtmp519 = in[946] & 1'b0;
	assign out[210] = in[1152] ^ in[137];
	assign out[246] = origtmp611 & in[57];
	assign origtmp1970 = origtmp2141 ^ origtmp1825;
	assign origtmp320 = origtmp318 | in[1268];
	assign out[185] = origtmp457 ^ origtmp458;
	assign origtmp342 = in[1073] | 1'b0;
	assign origtmp330 = 1'b0 & 1'b0;
	assign origtmp640 = ~in[364];
	assign origtmp594 = ~1'b1;
	assign origtmp1370 = in[1346] | in[321];
	assign origtmp487 = 1'b1 ^ 1'b1;
	assign origtmp1873 = in[1468] | in[515];
	assign origtmp1042 = origtmp1045 | 1'b0;
	assign origtmp17 = origtmp20 & origtmp20;
	assign origtmp281 = in[461] & in[461];
	assign origtmp1264 = in[1294] ^ origtmp1820;
	assign origtmp230 = ~origtmp231;
	assign origtmp2194 = in[288] ^ in[761];
	assign out[189] = origtmp470 | origtmp471;
	assign origtmp1265 = in[1337] ^ origtmp2081;
	assign out[54] = origtmp131;
	assign origtmp1949 = origtmp1479 | origtmp1812;
	assign origtmp1679 = origtmp1890 ^ origtmp2219;
	assign out[296] = origtmp746 & origtmp746;
	assign origtmp635 = in[368] | in[130];
	assign origtmp1822 = origtmp2056 ^ in[471];
	assign origtmp1230 = in[610] ^ origtmp1231;
	assign origtmp1184 = 1'b1 ^ 1'b1;
	assign origtmp1331 = in[763] | in[1369];
	assign origtmp305 = ~in[1439];
	assign origtmp515 = 1'b1;
	assign out[438] = 1'b1 & 1'b0;
	assign origtmp1716 = origtmp2164 & in[781];
	assign origtmp512 = origtmp513 | origtmp510;
	assign origtmp832 = 1'b0 ^ 1'b1;
	assign out[249] = in[1005] & origtmp620;
	assign out[120] = origtmp298 & origtmp297;
	assign origtmp2189 = origtmp1984 ^ in[147];
	assign origtmp1372 = in[753] ^ in[179];
	assign origtmp750 = 1'b1;
	assign origtmp360 = 1'b0 | in[1143];
	assign origtmp1308 = origtmp2151 & origtmp1829;
	assign out[405] = origtmp999 & in[602];
	assign origtmp1447 = origtmp1460 & in[1137];
	assign origtmp1149 = 1'b1 & in[653];
	assign origtmp924 = in[780] ^ in[116];
	assign origtmp739 = 1'b0 ^ origtmp737;
	assign origtmp816 = 1'b1 & origtmp818;
	assign origtmp1441 = origtmp1768 | origtmp2118;
	assign origtmp900 = origtmp901 & 1'b0;
	assign out[136] = origtmp335 ^ origtmp334;
	assign origtmp800 = in[1161] ^ 1'b1;
	assign out[155] = in[276] | 1'b0;
	assign origtmp1124 = in[273] & in[273];
	assign origtmp2138 = in[1397] ^ in[989];
	assign origtmp2090 = origtmp1932 ^ in[910];
	assign origtmp568 = origtmp571 ^ origtmp572;
	assign origtmp889 = in[2] & in[96];
	assign origtmp27 = ~1'b1;
	assign origtmp1934 = origtmp2211 & origtmp2229;
	assign origtmp538 = 1'b1 | origtmp539;
	assign origtmp1903 = in[734] ^ in[941];
	assign origtmp1448 = origtmp2206 ^ origtmp1502;
	assign origtmp329 = origtmp328 & in[146];
	assign origtmp1556 = in[84] | in[1119];
	assign origtmp1559 = origtmp1575 | in[217];
	assign origtmp1899 = origtmp2042 ^ origtmp1333;
	assign origtmp506 = 1'b1 & 1'b1;
	assign origtmp475 = in[738] | 1'b1;
	assign origtmp1260 = origtmp1743 | origtmp1894;
	assign origtmp763 = 1'b1 ^ in[695];
	assign origtmp557 = origtmp560 | 1'b0;
	assign origtmp1728 = in[497] | in[1088];
	assign origtmp2193 = in[1463] ^ in[434];
	assign origtmp1166 = in[787] | in[787];
	assign origtmp1568 = in[216] | in[419];
	assign origtmp18 = ~origtmp20;
	assign out[36] = origtmp96 & in[182];
	assign origtmp968 = origtmp971 & origtmp971;
	assign out[442] = in[898] | origtmp1097;
	assign origtmp1379 = origtmp1762 & origtmp2208;
	assign out[494] = origtmp1233 & in[627];
	assign origtmp770 = ~origtmp767;
	assign origtmp2176 = origtmp2139 ^ in[1224];
	assign origtmp2093 = in[448] | in[641];
	assign origtmp1294 = origtmp1270 ^ origtmp1422;
	assign origtmp1027 = in[1118] ^ 1'b0;
	assign origtmp176 = 1'b1 | 1'b1;
	assign origtmp2200 = origtmp1680 & in[1296];
	assign origtmp997 = 1'b1 & 1'b0;
	assign origtmp311 = 1'b1;
	assign origtmp2165 = in[81] ^ origtmp1283;
	assign origtmp405 = 1'b0 | 1'b1;
	assign origtmp1158 = 1'b0 ^ origtmp1157;
	assign origtmp1115 = origtmp1116 & 1'b1;
	assign origtmp1962 = in[868] | in[904];
	assign origtmp585 = in[519] | origtmp586;
	assign origtmp2149 = origtmp2049 | origtmp1840;
	assign out[202] = origtmp512 & in[1233];
	assign out[16] = origtmp38;
	assign origtmp1733 = in[405] | origtmp1551;
	assign origtmp1710 = origtmp1783 & in[601];
	assign origtmp708 = in[977] | in[1257];
	assign out[381] = origtmp938 | origtmp937;
	assign origtmp1320 = origtmp1557 ^ origtmp2230;
	assign origtmp661 = 1'b1 & 1'b0;
	assign origtmp1686 = in[1318] | in[895];
	assign origtmp1498 = origtmp2241 & origtmp2066;
	assign origtmp513 = origtmp511 ^ origtmp511;
	assign origtmp1 = in[544] | 1'b0;
	assign origtmp1298 = origtmp1997 | in[543];
	assign origtmp1770 = in[706] | origtmp1698;
	assign out[464] = origtmp1165 & 1'b1;
	assign origtmp720 = 1'b0 | 1'b0;
	assign origtmp1181 = ~in[1084];
	assign origtmp1891 = in[1177] | in[1027];
	assign origtmp1569 = origtmp1841 ^ origtmp1632;
	assign origtmp1723 = origtmp1411 | origtmp2204;
	assign origtmp2205 = origtmp1924 | origtmp1941;
	assign origtmp2002 = origtmp1332 ^ origtmp1329;
	assign origtmp263 = 1'b1 & origtmp264;
	assign origtmp530 = origtmp529 ^ in[1414];
	assign origtmp81 = 1'b0;
	assign out[425] = origtmp1055 | 1'b0;
	assign origtmp1036 = origtmp1035;
	assign origtmp2008 = origtmp1339 & in[219];
	assign origtmp1586 = in[839] & in[1392];
	assign origtmp1737 = in[578] | in[1455];
	assign origtmp1477 = origtmp1974 & origtmp1757;
	assign origtmp1756 = origtmp2169 ^ origtmp1980;
	assign origtmp1973 = in[1492] ^ in[344];
	assign origtmp1302 = in[1405] ^ origtmp1382;
	assign origtmp41 = ~origtmp39;
	assign origtmp601 = 1'b1 ^ 1'b0;
	assign origtmp660 = ~1'b0;
	assign origtmp132 = 1'b0 | in[1032];
	assign origtmp480 = origtmp477;
	assign origtmp798 = 1'b1 & in[1161];
	assign origtmp1164 = 1'b0 | 1'b0;
	assign origtmp1848 = origtmp1272 ^ origtmp2044;
	assign origtmp2029 = in[291] ^ in[705];
	assign origtmp954 = ~1'b1;
	assign origtmp1385 = origtmp1579 ^ in[1421];
	assign out[142] = origtmp353 ^ origtmp352;
	assign origtmp857 = origtmp856 & origtmp856;
	assign origtmp1330 = origtmp2064 & in[1225];
	assign origtmp870 = 1'b0 ^ 1'b0;
	assign origtmp266 = ~in[841];
	assign origtmp1145 = in[856];
	assign out[22] = origtmp55 ^ origtmp54;
	assign out[57] = origtmp140 | origtmp139;
	assign origtmp1495 = in[1090] | origtmp1242;
	assign origtmp2012 = origtmp2140 & in[438];
	assign origtmp196 = 1'b1 | in[91];
	assign out[158] = in[545] ^ in[340];
	assign origtmp1489 = origtmp1559 | in[423];
	assign origtmp1263 = in[806] & origtmp1790;
	assign origtmp598 = ~1'b0;
	assign origtmp1598 = origtmp1492 & origtmp1961;
	assign origtmp1900 = in[490] ^ origtmp1374;
	assign out[60] = origtmp148 | origtmp147;
	assign origtmp707 = 1'b0 | origtmp704;
	assign origtmp648 = origtmp649 ^ origtmp646;
	assign out[145] = origtmp359 ^ in[420];
	assign origtmp2146 = origtmp1518 & origtmp1495;
	assign origtmp804 = in[1226] ^ in[1226];
	assign origtmp280 = 1'b0;
	assign origtmp1642 = origtmp1486 ^ origtmp1765;
	assign origtmp623 = 1'b0;
	assign origtmp2119 = origtmp1271 ^ in[526];
	assign origtmp309 = 1'b0;
	assign origtmp2254 = origtmp1970 & origtmp1315;
	assign origtmp1959 = origtmp2120 & in[459];
	assign origtmp1578 = origtmp1816 | origtmp1674;
	assign origtmp1984 = in[1046] | in[552];
	assign out[419] = origtmp1033 ^ origtmp1031;
	assign origtmp787 = ~origtmp788;
	assign origtmp1786 = origtmp1740 & in[38];
	assign origtmp43 = 1'b0 | 1'b0;
	assign origtmp1874 = origtmp1718 | origtmp1250;
	assign origtmp1538 = origtmp1365 | origtmp1838;
	assign origtmp2067 = origtmp1477 & origtmp1712;
	assign out[351] = origtmp875 & origtmp876;
	assign origtmp689 = origtmp687 & origtmp688;
	assign origtmp1799 = in[174] ^ in[1232];
	assign origtmp543 = 1'b1;
	assign origtmp1352 = origtmp2131 | origtmp1581;
	assign origtmp1059 = 1'b1;
	assign origtmp1281 = origtmp1802 & in[1210];
	assign origtmp932 = 1'b0 & in[719];
	assign origtmp292 = in[537] & in[1164];
	assign out[154] = origtmp383;
	assign origtmp2088 = origtmp1865 | origtmp1278;
	assign origtmp833 = ~origtmp832;
	assign out[263] = 1'b1 ^ origtmp650;
	assign out[175] = in[606] ^ origtmp440;
	assign origtmp326 = in[146] & 1'b1;
	assign origtmp87 = 1'b1 | 1'b0;
	assign origtmp1130 = 1'b1 & 1'b0;
	assign origtmp504 = in[822] | 1'b0;
	assign origtmp1187 = 1'b0 | 1'b1;
	assign origtmp1173 = ~in[1246];
	assign origtmp2237 = in[889] ^ origtmp2039;
	assign origtmp2007 = origtmp1543 | origtmp1830;
	assign origtmp806 = in[464] ^ in[492];
	assign origtmp1396 = origtmp1655 ^ in[117];
	assign origtmp1842 = origtmp2037 & in[727];
	assign origtmp877 = in[1395] | in[1395];
	assign origtmp508 = origtmp506 | origtmp509;
	assign origtmp1258 = in[232] | in[1222];
	assign origtmp1051 = origtmp1048 ^ origtmp1048;
	assign origtmp1815 = origtmp2225 | origtmp1352;
	assign origtmp2064 = in[263] | in[186];
	assign origtmp1351 = in[881] & in[848];
	assign origtmp1161 = in[13] & origtmp1159;
	assign origtmp335 = in[1323] | in[852];
	assign origtmp378 = ~1'b1;
	assign out[198] = origtmp498;
	assign origtmp170 = 1'b1;
	assign origtmp234 = origtmp230 ^ 1'b1;
	assign out[315] = in[1489] & in[55];
	assign out[197] = origtmp497 | origtmp495;
	assign origtmp377 = ~1'b1;
	assign origtmp592 = origtmp594 & origtmp594;
	assign origtmp957 = origtmp956 ^ in[672];
	assign origtmp135 = origtmp132 | origtmp133;
	assign out[149] = origtmp371 & origtmp367;
	assign origtmp1536 = in[337] | in[1049];
	assign origtmp980 = origtmp981 ^ origtmp981;
	assign origtmp1774 = origtmp2033 ^ in[160];
	assign origtmp1082 = 1'b0 ^ 1'b1;
	assign origtmp1162 = ~1'b1;
	assign origtmp2139 = in[1191] | origtmp1494;
	assign origtmp974 = ~in[536];
	assign origtmp1706 = origtmp1525 | origtmp1299;
	assign origtmp569 = in[520] & 1'b0;
	assign origtmp2010 = origtmp2210 ^ origtmp1887;
	assign origtmp978 = 1'b0 & 1'b1;
	assign origtmp413 = in[443] & 1'b1;
	assign out[13] = 1'b0 ^ 1'b0;
	assign origtmp1193 = origtmp1192 ^ 1'b1;
	assign origtmp7 = 1'b0 ^ in[634];
	assign origtmp1868 = origtmp1681 | in[1108];
	assign origtmp1721 = in[1467] ^ in[576];
	assign origtmp2126 = in[249] ^ in[548];
	assign origtmp2109 = origtmp1542 ^ origtmp1785;
	assign origtmp1493 = origtmp2087 & origtmp1990;
	assign origtmp341 = 1'b0 & 1'b1;
	assign origtmp186 = origtmp185 ^ origtmp185;
	assign origtmp675 = 1'b1 | origtmp674;
	assign origtmp110 = 1'b1;
	assign origtmp1101 = 1'b0;
	assign origtmp1615 = in[599] ^ origtmp1753;
	assign out[290] = ~in[1227];
	assign origtmp129 = 1'b1 & in[1097];
	assign out[2] = origtmp4 & origtmp5;
	assign out[318] = ~1'b0;
	assign origtmp1834 = in[643] | origtmp1751;
	assign origtmp228 = 1'b0 ^ in[676];
	assign origtmp454 = 1'b1 & origtmp453;
	assign origtmp1432 = in[367] | in[1069];
	assign origtmp94 = origtmp93 & in[796];
	assign out[9] = origtmp21 | origtmp19;
	assign out[370] = origtmp911 | origtmp910;
	assign origtmp646 = 1'b1 & origtmp647;
	assign origtmp1846 = origtmp1620 | in[1424];
	assign origtmp1795 = origtmp1497 | origtmp1835;
	assign out[123] = origtmp304 & 1'b0;
	assign origtmp1935 = in[1319] ^ origtmp1982;
	assign origtmp383 = origtmp385 | in[384];
	assign origtmp801 = origtmp800 & in[747];
	assign origtmp1892 = origtmp1421 & origtmp2027;
	assign out[423] = origtmp1047 | origtmp1046;
	assign origtmp1267 = in[264] | origtmp1899;
	assign origtmp2188 = in[283] ^ origtmp1531;
	assign origtmp1160 = ~origtmp1161;
	assign origtmp1885 = origtmp1993 & origtmp2181;
	assign origtmp218 = 1'b0 | origtmp217;
	assign origtmp1484 = in[400] & in[1478];
	assign origtmp306 = origtmp308 ^ in[1439];
	assign origtmp1033 = 1'b0 & origtmp1032;
	assign origtmp1024 = 1'b1 ^ 1'b1;
	assign origtmp784 = origtmp785 & origtmp785;
	assign origtmp262 = ~1'b0;
	assign origtmp852 = in[1250] & in[1250];
	assign origtmp84 = origtmp85 & in[123];
	assign origtmp1628 = in[523] ^ in[1012];
	assign origtmp2221 = in[1390] & in[668];
	assign origtmp831 = origtmp832 & 1'b1;
	assign origtmp1313 = origtmp2021 & origtmp2238;
	assign origtmp651 = 1'b1;
	assign origtmp703 = origtmp702;
	assign origtmp789 = origtmp791 | origtmp790;
	assign origtmp232 = origtmp231 & origtmp231;
	assign origtmp1636 = in[52] | in[785];
	assign origtmp993 = 1'b1 & in[1020];
	assign origtmp890 = in[1229] | in[120];
	assign origtmp2078 = in[1194] ^ origtmp1370;
	assign origtmp735 = in[767] & 1'b1;
	assign origtmp1012 = 1'b0 & in[24];
	assign origtmp525 = in[891] | in[422];
	assign origtmp1156 = 1'b0;
	assign origtmp2066 = origtmp1515 | origtmp1707;
	assign origtmp671 = origtmp673 ^ in[1100];
	assign origtmp1222 = 1'b0 ^ in[708];
	assign out[369] = 1'b1 ^ origtmp909;
	assign out[427] = origtmp1062 & origtmp1063;
	assign origtmp1877 = origtmp2108 | in[331];
	assign origtmp1407 = origtmp1621 & in[966];
	assign origtmp1252 = in[964] ^ in[654];
	assign origtmp49 = in[905] & origtmp50;
	assign origtmp2203 = in[663] & origtmp1807;
	assign origtmp1555 = origtmp1747 & origtmp1400;
	assign origtmp1796 = in[1110] & in[1016];
	assign origtmp106 = ~in[496];
	assign out[424] = origtmp1051 | 1'b1;
	assign origtmp237 = 1'b1 ^ 1'b0;
	assign origtmp382 = in[124] ^ in[1315];
	assign origtmp1813 = origtmp1325 & origtmp1395;
	assign origtmp1597 = in[901] | in[795];
	assign origtmp2145 = origtmp1898 | origtmp1457;
	assign origtmp2127 = in[435] & in[272];
	assign out[98] = in[585] & in[585];
	assign origtmp1405 = origtmp1949 & origtmp1553;
	assign origtmp559 = 1'b1 ^ 1'b0;
	assign origtmp344 = in[228] ^ origtmp347;
	assign origtmp1132 = in[818] & in[90];
	assign out[373] = origtmp921 & origtmp920;
	assign origtmp1099 = origtmp1100 | in[1258];
	assign origtmp1009 = origtmp1008;
	assign out[30] = in[1139] | 1'b0;
	assign origtmp755 = in[1331] | origtmp756;
	assign out[420] = 1'b0 | origtmp1037;
	assign origtmp148 = 1'b1 ^ in[241];
	assign origtmp1153 = 1'b1 ^ origtmp1152;
	assign origtmp1073 = 1'b0 & 1'b1;
	assign out[303] = origtmp760 ^ 1'b1;
	assign origtmp926 = in[478] & in[354];
	assign origtmp351 = 1'b0 | 1'b1;
	assign origtmp1768 = origtmp2213 | origtmp1704;
	assign origtmp951 = 1'b1;
	assign out[208] = 1'b0 | origtmp516;
	assign origtmp1777 = in[385] & in[1349];
	assign origtmp439 = origtmp438 ^ origtmp438;
	assign out[29] = 1'b1 | origtmp78;
	assign origtmp387 = 1'b0;
	assign origtmp1798 = origtmp2135 | origtmp1440;
	assign origtmp202 = ~origtmp204;
	assign origtmp1695 = origtmp1509 | origtmp1429;
	assign origtmp2153 = in[1291] | origtmp1574;
	assign out[201] = origtmp508 & origtmp507;
	assign origtmp656 = ~origtmp655;
	assign origtmp1072 = 1'b0 | origtmp1070;
	assign origtmp1290 = origtmp2032 & origtmp1343;
	assign out[69] = 1'b1 ^ in[166];
	assign origtmp52 = in[513] | 1'b1;
	assign origtmp29 = ~1'b0;
	assign origtmp827 = origtmp826 | in[1458];
	assign origtmp1787 = in[678] ^ in[1300];
	assign origtmp1328 = origtmp1368 | origtmp1301;
	assign origtmp239 = in[1293];
	assign origtmp1691 = in[51] ^ in[247];
	assign origtmp575 = in[417] & in[315];
	assign out[417] = in[1289] ^ origtmp1026;
	assign origtmp2048 = in[149] | in[173];
	assign origtmp373 = origtmp376;
	assign origtmp1582 = in[356] | in[1360];
	assign origtmp1930 = origtmp1424 | origtmp2199;
	assign origtmp945 = origtmp946 ^ in[1350];
	assign origtmp287 = 1'b0;
	assign out[188] = origtmp466 & origtmp466;
	assign origtmp1109 = in[505];
	assign origtmp1431 = in[859] ^ origtmp2119;
	assign origtmp1389 = in[742] | origtmp1412;
	assign origtmp2201 = in[407] | in[86];
	assign origtmp83 = in[123];
	assign origtmp2181 = in[1011] | in[415];
	assign origtmp1592 = origtmp1324 ^ in[1215];
	assign origtmp955 = 1'b1 & origtmp952;
	assign origtmp1859 = origtmp1556 ^ origtmp1985;
	assign origtmp138 = origtmp137 & in[843];
	assign origtmp642 = 1'b0 | origtmp641;
	assign origtmp2037 = in[17] | origtmp1398;
	assign origtmp567 = in[99] ^ 1'b1;
	assign out[451] = origtmp1128;
	assign origtmp1793 = origtmp1408 | origtmp2022;
	assign origtmp2009 = in[1180] | in[305];
	assign origtmp187 = origtmp186;
	assign origtmp1400 = in[579] | in[336];
	assign origtmp1044 = origtmp1042 & origtmp1042;
	assign out[85] = origtmp209 ^ origtmp209;
	assign origtmp1806 = in[1333] ^ in[624];
	assign origtmp255 = ~in[112];
	assign out[432] = 1'b1 | origtmp1073;
	assign out[260] = origtmp644 | 1'b0;
	assign origtmp251 = origtmp252 & origtmp252;
	assign origtmp1674 = origtmp1501 & origtmp1461;
	assign origtmp563 = 1'b0 & 1'b0;
	assign origtmp1740 = in[1037] | in[598];
	assign origtmp1217 = in[1412] & in[1412];
	assign out[4] = in[735] & in[1344];
	assign origtmp1760 = in[1038] ^ in[907];
	assign origtmp670 = ~in[1100];
	assign origtmp257 = in[670] & origtmp260;
	assign origtmp12 = 1'b0 | 1'b1;
	assign origtmp1089 = 1'b0 | origtmp1091;
	assign origtmp753 = origtmp752;
	assign origtmp447 = in[1197] ^ in[1197];
	assign origtmp915 = in[1098] & in[1098];
	assign origtmp67 = in[952] & origtmp66;
	assign origtmp746 = in[1329];
	assign out[240] = in[595] | origtmp599;
	assign origtmp2255 = in[764] | origtmp1425;
	assign origtmp1362 = origtmp1773 ^ origtmp1973;
	assign out[50] = origtmp124 | origtmp123;
	assign origtmp1784 = in[1156] | origtmp1957;
	assign out[147] = origtmp363 & origtmp364;
	assign out[437] = origtmp1085 ^ origtmp1085;
	assign origtmp1932 = in[662] & in[1025];
	assign out[94] = in[1357] | origtmp235;
	assign origtmp1131 = origtmp1133 | in[90];
	assign origtmp943 = 1'b1;
	assign origtmp1986 = origtmp1441 ^ origtmp1584;
	assign origtmp673 = in[1100] ^ in[162];
	assign out[334] = origtmp836 ^ origtmp834;
	assign origtmp984 = origtmp983 & origtmp982;
	assign origtmp10 = in[1474] ^ origtmp9;
	assign out[34] = ~origtmp92;
	assign origtmp1199 = origtmp1196 | origtmp1195;
	assign out[258] = origtmp643 | origtmp642;
	assign out[259] = in[1495] | in[1345];
	assign out[70] = in[984] & 1'b0;
	assign out[288] = origtmp729 | 1'b0;
	assign origtmp2225 = in[739] ^ in[791];
	assign origtmp1808 = in[204] | in[532];
	assign origtmp1727 = origtmp1701 | origtmp1880;
	assign origtmp1722 = origtmp2090 | origtmp2077;
	assign origtmp1361 = origtmp1583 | origtmp1562;
	assign origtmp2163 = origtmp2178 & in[1162];
	assign origtmp1271 = origtmp1321 | in[144];
	assign origtmp225 = in[960];
	assign origtmp1888 = origtmp2156 ^ origtmp1643;
	assign origtmp878 = in[1010] & origtmp880;
	assign origtmp873 = origtmp872 & origtmp872;
	assign origtmp658 = in[431] & 1'b1;
	assign out[216] = origtmp533 & origtmp536;
	assign origtmp1961 = origtmp1393 | in[718];
	assign origtmp1227 = origtmp1228 | origtmp1225;
	assign origtmp1705 = origtmp1251 ^ origtmp1407;
	assign origtmp402 = origtmp399 & origtmp400;
	assign origtmp1421 = in[605] ^ origtmp1356;
	assign origtmp1711 = origtmp2255 ^ origtmp1453;
	assign origtmp371 = ~origtmp370;
	assign origtmp1832 = in[94] | in[940];
	assign origtmp1047 = in[816] | 1'b0;
	assign out[403] = in[1064];
	assign origtmp1434 = origtmp1842 | in[18];
	assign out[17] = origtmp39 ^ origtmp41;
	assign origtmp1107 = origtmp1108 | origtmp1106;
	assign out[257] = 1'b1 ^ origtmp637;
	assign origtmp1526 = origtmp2149 | origtmp2099;
	assign origtmp1338 = in[1150] ^ origtmp1532;
	assign out[407] = origtmp1002;
	assign origtmp1678 = origtmp1647 & origtmp1630;
	assign origtmp1714 = in[916] & in[67];
	assign origtmp571 = in[520] ^ in[520];
	assign origtmp1872 = in[408] & origtmp1749;
	assign origtmp906 = ~1'b1;
	assign origtmp2180 = in[1124] ^ origtmp2115;
	assign origtmp1225 = in[79] & in[79];
	assign origtmp987 = in[163] & 1'b0;
	assign origtmp916 = in[168] | 1'b1;
	assign origtmp652 = origtmp651;
	assign origtmp649 = 1'b0 & origtmp647;
	assign origtmp425 = origtmp424 & 1'b1;
	assign origtmp1127 = origtmp1126 | in[1216];
	assign out[53] = in[106] & in[374];
	assign origtmp1046 = 1'b0 ^ in[816];
	assign origtmp397 = origtmp396 | origtmp396;
	assign origtmp209 = origtmp210 | origtmp208;
	assign out[485] = in[338] ^ in[1339];
	assign out[14] = origtmp31 | origtmp29;
	assign origtmp443 = origtmp444 ^ 1'b1;
	assign origtmp1104 = origtmp1101 & origtmp1102;
	assign origtmp380 = in[1315] & origtmp381;
	assign origtmp1038 = 1'b1 & 1'b1;
	assign origtmp562 = origtmp566 | origtmp563;
	assign origtmp696 = origtmp697 | origtmp697;
	assign origtmp884 = in[297] | origtmp883;
	assign origtmp2208 = origtmp1289 | origtmp1875;
	assign origtmp92 = origtmp91 ^ origtmp94;
	assign origtmp1850 = origtmp1406 & origtmp1304;
	assign origtmp785 = ~1'b0;
	assign origtmp863 = origtmp864 & origtmp865;
	assign origtmp2171 = origtmp1981 & in[440];
	assign out[200] = origtmp505 & origtmp504;
	assign out[307] = in[1435] | in[1230];
	assign origtmp1341 = in[1267] | in[260];
	assign origtmp1087 = 1'b1 & origtmp1088;
	assign out[489] = ~1'b1;
	assign origtmp1996 = in[522] & in[1198];
	assign origtmp2169 = in[893] & origtmp1437;
	assign origtmp1902 = origtmp2142 & origtmp1318;
	assign out[243] = origtmp606 & origtmp605;
	assign origtmp861 = 1'b0 | origtmp859;
	assign origtmp96 = 1'b0 | 1'b0;
	assign origtmp254 = origtmp255 & 1'b0;
	assign origtmp2084 = origtmp2123 ^ origtmp1597;
	assign origtmp2168 = in[924] ^ in[319];
	assign origtmp278 = 1'b0 | 1'b0;
	assign origtmp1931 = in[329] | origtmp1789;
	assign out[8] = origtmp14 ^ origtmp15;
	assign origtmp1647 = in[529] | origtmp1937;
	assign origtmp1968 = in[880] & in[617];
	assign out[346] = origtmp861 & origtmp862;
	assign origtmp1392 = origtmp2159 & origtmp1611;
	assign origtmp107 = 1'b0 ^ in[496];
	assign origtmp1134 = origtmp1135 & origtmp1135;
	assign origtmp553 = in[479] & origtmp554;
	assign origtmp663 = origtmp661 ^ 1'b1;
	assign origtmp1571 = origtmp1615 & in[983];
	assign origtmp1188 = 1'b0 | 1'b0;
	assign origtmp1103 = ~origtmp1104;
	assign out[187] = origtmp463 & in[842];
	assign origtmp1522 = in[1422] ^ origtmp1607;
	assign origtmp1866 = in[618] | in[1427];
	assign origtmp1068 = origtmp1071 & 1'b0;
	assign origtmp2019 = origtmp1994 ^ origtmp1526;
	assign origtmp769 = 1'b0 ^ in[884];
	assign origtmp2015 = in[1114] & in[1490];
	assign origtmp1993 = origtmp2023 ^ in[277];
	assign origtmp1880 = origtmp1792 | in[1407];
	assign origtmp1088 = 1'b0;
	assign out[306] = origtmp768 | origtmp770;
	assign out[184] = 1'b1 & origtmp454;
	assign origtmp22 = 1'b0 | 1'b0;
	assign origtmp466 = 1'b1 & origtmp467;
	assign origtmp1002 = origtmp1001 ^ 1'b1;
	assign origtmp1958 = origtmp1808 & in[1321];
	assign origtmp363 = 1'b0 & origtmp365;
	assign origtmp872 = 1'b0;
	assign origtmp245 = 1'b1 & 1'b0;
	assign origtmp1311 = in[1072] ^ in[571];
	assign origtmp364 = 1'b0 ^ 1'b1;
	assign out[194] = ~in[892];
	assign origtmp1606 = in[788] ^ origtmp2240;
	assign out[164] = origtmp410 | 1'b0;
	assign origtmp422 = 1'b1;
	assign origtmp2234 = in[475] & origtmp2105;
	assign origtmp786 = origtmp785;
	assign origtmp412 = in[949] & in[1094];
	assign out[324] = in[492] & origtmp806;
	assign origtmp1118 = origtmp1116 ^ in[541];
	assign origtmp130 = in[642] ^ in[642];
	assign origtmp888 = 1'b0;
	assign origtmp551 = 1'b1 | in[721];
	assign origtmp2198 = origtmp1652 & origtmp1794;
	assign origtmp61 = origtmp63 | in[189];
	assign out[426] = origtmp1060 ^ origtmp1057;
	assign origtmp1844 = in[982] & in[652];
	assign origtmp518 = origtmp519 ^ 1'b1;
	assign origtmp144 = in[1336] | in[1336];
	assign out[453] = origtmp1131 ^ origtmp1132;
	assign out[353] = origtmp879 & origtmp881;
	assign origtmp2027 = in[883] ^ in[584];
	assign origtmp1707 = in[183] ^ origtmp1414;
	assign out[65] = origtmp165 ^ origtmp167;
	assign origtmp1637 = in[962] ^ in[798];
	assign origtmp166 = origtmp164 ^ origtmp164;
	assign out[492] = origtmp1227 ^ origtmp1229;
	assign origtmp1345 = origtmp1466 | in[493];
	assign origtmp1186 = origtmp1185 & origtmp1183;
	assign out[274] = ~origtmp689;
	assign origtmp1496 = origtmp1292 | origtmp1381;
	assign origtmp435 = origtmp434 | origtmp432;
	assign origtmp2191 = in[1057] | origtmp2114;
	assign origtmp1097 = in[582] ^ 1'b1;
	assign out[151] = origtmp379 ^ origtmp378;
	assign origtmp981 = ~in[463];
	assign origtmp759 = 1'b0;
	assign origtmp1546 = origtmp1371 & origtmp1695;
	assign origtmp1861 = in[975] | in[945];
	assign origtmp1077 = in[1309] & origtmp1074;
	assign origtmp112 = in[1416] & in[1416];
	assign origtmp1071 = 1'b0;
	assign origtmp246 = 1'b0;
	assign origtmp1830 = origtmp2144 & in[1113];
	assign origtmp2174 = origtmp1796 ^ origtmp1350;
	assign origtmp2065 = in[1342] ^ in[1023];
	assign origtmp1732 = origtmp2083 & origtmp2184;
	assign origtmp782 = in[502] & 1'b0;
	assign origtmp346 = origtmp345 ^ origtmp343;
	assign origtmp80 = origtmp81 ^ origtmp77;
	assign origtmp114 = origtmp113 | in[701];
	assign origtmp1223 = origtmp1220 | 1'b1;
	assign origtmp2152 = in[78] | origtmp2053;
	assign origtmp741 = origtmp740;
	assign origtmp250 = 1'b0 & 1'b1;
	assign origtmp511 = in[1233] ^ 1'b0;
	assign origtmp161 = 1'b1 | in[360];
	assign origtmp2018 = origtmp1379 | in[317];
	assign origtmp1272 = origtmp1567 | in[41];
	assign out[66] = origtmp169 ^ origtmp169;
	assign out[141] = 1'b0 ^ origtmp348;
	assign out[379] = in[436] | 1'b0;
	assign out[47] = origtmp114 | origtmp113;
	assign origtmp1682 = origtmp2024 | in[129];
	assign out[131] = 1'b0 ^ 1'b0;
	assign origtmp865 = 1'b1 ^ in[148];
	assign origtmp1651 = in[756] & in[1213];
	assign origtmp956 = 1'b0 | in[672];
	assign origtmp774 = origtmp772;
	assign origtmp160 = 1'b0 & origtmp161;
	assign out[169] = origtmp419 ^ origtmp420;
	assign out[238] = origtmp590 ^ origtmp591;
	assign origtmp24 = 1'b0 | origtmp26;
	assign origtmp1032 = in[1123] & origtmp1034;
	assign origtmp1159 = origtmp1158 & in[13];
	assign origtmp1070 = origtmp1069 ^ origtmp1068;
	assign origtmp1137 = in[1383] ^ 1'b1;
	assign origtmp2030 = in[1340] | origtmp1983;
	assign origtmp2247 = in[239] & in[1081];
	assign out[280] = origtmp706 ^ origtmp707;
	assign origtmp637 = origtmp639 ^ origtmp638;
	assign out[261] = origtmp648;
	assign origtmp970 = origtmp968 | origtmp972;
	assign origtmp2120 = origtmp1560 | in[445];
	assign origtmp1343 = origtmp2094 ^ origtmp1341;
	assign origtmp862 = origtmp860 & in[138];
	assign origtmp958 = origtmp959 & origtmp957;
	assign origtmp1163 = 1'b0 | origtmp1162;
	assign origtmp547 = 1'b1;
	assign origtmp284 = origtmp285;
	assign out[327] = origtmp813 & 1'b1;
	assign origtmp1102 = ~in[1047];
	assign origtmp1790 = origtmp2126 & in[85];
	assign out[414] = origtmp1018 ^ origtmp1020;
	assign origtmp1769 = in[849] & in[1461];
	assign origtmp1490 = in[218] ^ in[1358];
	assign origtmp1414 = in[229] | in[1208];
	assign origtmp1209 = 1'b1 | 1'b1;
	assign origtmp666 = 1'b1;
	assign origtmp1627 = in[1260] ^ in[675];
	assign origtmp1667 = origtmp1416 & origtmp1815;
	assign origtmp843 = in[640];
	assign out[83] = 1'b0 ^ 1'b0;
	assign origtmp1471 = origtmp1439 ^ origtmp1905;
	assign origtmp103 = in[504] | origtmp101;
	assign origtmp496 = 1'b0;
	assign origtmp446 = 1'b1 & 1'b0;
	assign out[21] = in[817] & in[817];
	assign origtmp722 = ~1'b0;
	assign origtmp1776 = origtmp2018 ^ origtmp1971;
	assign origtmp1755 = in[205] | in[547];
	assign out[37] = origtmp98 ^ origtmp98;
	assign origtmp1901 = origtmp1956 ^ origtmp2055;
	assign origtmp626 = 1'b1;
	assign origtmp211 = 1'b1 ^ 1'b0;
	assign origtmp1458 = in[233] ^ in[382];
	assign origtmp1766 = in[1449] | in[648];
	assign origtmp983 = in[1253] | origtmp986;
	assign origtmp1170 = origtmp1172;
	assign origtmp2036 = in[93] | origtmp1402;
	assign origtmp312 = origtmp313 | origtmp311;
	assign origtmp159 = origtmp157;
	assign origtmp2155 = in[5] | in[1201];
	assign out[1] = origtmp2 | 1'b1;
	assign origtmp1574 = in[396] | origtmp2059;
	assign origtmp1539 = in[1183] & in[342];
	assign origtmp1045 = 1'b0 ^ 1'b0;
	assign origtmp710 = in[697] | origtmp711;
	assign origtmp1856 = in[725] | in[199];
	assign origtmp2244 = in[1374] ^ in[290];
	assign origtmp25 = ~1'b0;
	assign origtmp1017 = 1'b0 ^ 1'b1;
	assign origtmp549 = origtmp548 ^ in[721];
	assign out[133] = origtmp329 & origtmp327;
	assign origtmp2059 = in[1131] | in[777];
	assign origtmp1524 = in[1103] & in[677];
	assign origtmp1394 = in[629] ^ in[6];
	assign origtmp1839 = in[421] | in[19];
	assign origtmp8 = origtmp7 ^ in[1486];
	assign origtmp768 = in[884] ^ in[884];
	assign origtmp350 = in[1004] & in[1004];
	assign origtmp1025 = 1'b1 ^ origtmp1024;
	assign origtmp841 = 1'b1;
	assign origtmp1952 = in[597] & in[1092];
	assign out[408] = origtmp1003 | 1'b0;
	assign origtmp1554 = in[326] & origtmp1967;
	assign out[433] = origtmp1076 & origtmp1077;
	assign origtmp866 = origtmp864 ^ origtmp863;
	assign out[51] = origtmp128 ^ origtmp127;
	assign origtmp1849 = origtmp1670 | origtmp1295;
	assign origtmp613 = origtmp615 ^ origtmp612;
	assign origtmp1907 = origtmp1864 & in[814];
	assign origtmp1611 = in[153] & origtmp1277;
	assign out[305] = in[784] ^ origtmp765;
	assign origtmp1413 = in[1217] & in[56];
	assign origtmp2157 = origtmp1569 | origtmp1929;
	assign origtmp2117 = origtmp1800 ^ origtmp1928;
	assign origtmp1869 = in[783] & in[1080];
	assign origtmp634 = origtmp635 ^ in[368];
	assign origtmp2150 = origtmp1510 | origtmp2254;
	assign origtmp1461 = origtmp2146 ^ origtmp1386;
	assign origtmp1356 = in[457] ^ in[1494];
	assign out[393] = origtmp973 | origtmp976;
	assign origtmp301 = origtmp302 & origtmp299;
	assign origtmp1912 = in[1207] & in[1354];
	assign origtmp630 = in[1460] | 1'b1;
	assign origtmp1879 = in[1359] & in[538];
	assign origtmp498 = in[256] & in[256];
	assign origtmp935 = in[719] ^ 1'b0;
	assign origtmp169 = 1'b0 | origtmp168;
	assign origtmp907 = 1'b1 & 1'b0;
	assign origtmp158 = origtmp157 | origtmp159;
	assign origtmp1506 = in[150] ^ in[717];
	assign origtmp1454 = in[1242] ^ in[267];
	assign origtmp855 = 1'b1 | 1'b1;
	assign origtmp90 = origtmp88 | origtmp89;
	assign origtmp1393 = origtmp2247 | origtmp1770;
	assign origtmp869 = in[70];
	assign out[449] = origtmp1119 | origtmp1117;
	assign origtmp1291 = origtmp1449 & origtmp1725;
	assign origtmp416 = in[510] ^ origtmp415;
	assign origtmp922 = in[361] & in[361];
	assign origtmp665 = 1'b0 & in[633];
	assign origtmp1587 = in[827] | in[1324];
	assign origtmp1108 = 1'b1 | 1'b1;
	assign origtmp1563 = in[703] | in[348];
	assign origtmp539 = ~origtmp537;
	assign origtmp657 = 1'b1 & 1'b0;
	assign origtmp1527 = in[728] & in[1052];
	assign origtmp126 = origtmp125 | in[430];
	assign origtmp481 = 1'b0;
	assign origtmp13 = origtmp16 & 1'b1;
	assign origtmp1701 = in[1041] | in[1306];
	assign origtmp1312 = origtmp1530 & origtmp1438;
	assign origtmp1235 = 1'b0 | 1'b0;
	assign out[241] = ~in[1393];
	assign out[125] = origtmp317 | origtmp316;
	assign out[264] = origtmp654 | origtmp657;
	assign origtmp795 = ~1'b1;
	assign origtmp937 = origtmp940 ^ origtmp939;
	assign origtmp1600 = origtmp1781 & origtmp1963;
	assign origtmp767 = origtmp771 | 1'b0;
	assign origtmp2042 = origtmp1940 & in[572];
	assign out[446] = 1'b0 ^ 1'b0;
	assign out[374] = ~1'b1;
	assign origtmp1745 = origtmp2129 | origtmp1622;
	assign origtmp830 = 1'b1 & 1'b0;
	assign origtmp1741 = in[107] | in[740];
	assign origtmp1964 = origtmp1741 & in[1054];
	assign out[182] = origtmp451 ^ origtmp449;
	assign out[447] = ~origtmp1110;
	assign origtmp418 = origtmp417 ^ in[255];
	assign origtmp2051 = in[1376] ^ in[1473];
	assign origtmp1649 = origtmp1760 & origtmp1505;
	assign origtmp1114 = origtmp1112 ^ 1'b1;
	assign origtmp1106 = origtmp1109 ^ origtmp1109;
	assign origtmp989 = in[412];
	assign origtmp1988 = origtmp1328 | origtmp1870;
	assign out[474] = 1'b1 | 1'b1;
	assign origtmp389 = ~in[9];
	assign origtmp1422 = in[900] & origtmp1446;
	assign origtmp517 = in[946] | origtmp518;
	assign origtmp2184 = in[140] ^ in[1484];
	assign origtmp1549 = in[26] ^ in[295];
	assign origtmp1232 = origtmp1230 & 1'b0;
	assign origtmp874 = ~1'b1;
	assign origtmp913 = ~origtmp915;
	assign out[58] = in[1051] & origtmp141;
	assign origtmp1327 = origtmp2045 | origtmp1496;
	assign origtmp1818 = in[956] ^ origtmp1305;
	assign out[62] = origtmp156 | 1'b1;
	assign origtmp1617 = origtmp1420 | origtmp1968;
	assign origtmp992 = ~origtmp991;
	assign origtmp1154 = origtmp1155 | origtmp1152;
	assign out[93] = origtmp234 | origtmp233;
	assign origtmp2099 = origtmp2127 | origtmp2034;
	assign origtmp1577 = origtmp2203 | in[418];
	assign origtmp182 = 1'b0 ^ 1'b0;
	assign origtmp1911 = in[923] ^ origtmp1799;
	assign origtmp71 = 1'b1 & 1'b0;
	assign origtmp490 = 1'b1;
	assign origtmp1533 = in[1175] ^ in[803];
	assign out[172] = in[82] & in[751];
	assign origtmp2161 = in[1158] | in[1436];
	assign origtmp2213 = origtmp2071 & origtmp2010;
	assign origtmp395 = origtmp392 & origtmp393;
	assign origtmp778 = origtmp775 ^ origtmp777;
	assign out[465] = origtmp1167 & origtmp1166;
	assign origtmp1835 = in[69] & in[355];
	assign origtmp736 = in[500] ^ origtmp738;
	assign origtmp2215 = origtmp1290 ^ origtmp1418;
	assign origtmp688 = 1'b0 & 1'b1;
	assign origtmp2058 = origtmp1244 | origtmp2111;
	assign origtmp1783 = origtmp1934 ^ origtmp1298;
	assign origtmp1929 = in[857] & origtmp1989;
	assign origtmp691 = origtmp692 ^ 1'b1;
	assign origtmp1491 = origtmp1297 & in[1347];
	assign origtmp247 = in[346] & in[346];
	assign origtmp1244 = in[1075] ^ in[1059];
	assign origtmp494 = origtmp491 ^ origtmp491;
	assign origtmp2044 = origtmp1264 & origtmp1570;
	assign origtmp609 = 1'b1;
	assign out[105] = origtmp261 | origtmp263;
	assign origtmp1023 = origtmp1024;
	assign origtmp1829 = origtmp2035 ^ origtmp1933;
	assign origtmp1376 = in[462] ^ origtmp1384;
	assign origtmp1395 = in[1425] | origtmp1541;
	assign out[90] = origtmp226 ^ origtmp225;
	assign origtmp2162 = origtmp2068 | in[132];
	assign origtmp552 = ~1'b0;
	assign origtmp599 = 1'b0 ^ origtmp598;
	assign origtmp886 = 1'b0 ^ 1'b1;
	assign origtmp880 = in[1010] & in[1010];
	assign out[301] = origtmp757 | origtmp758;
	assign origtmp1983 = origtmp2106 ^ origtmp2239;
	assign origtmp677 = 1'b1 | in[1067];
	assign origtmp69 = origtmp71 ^ 1'b1;
	assign origtmp274 = 1'b0 | 1'b0;
	assign origtmp1653 = in[837] ^ origtmp1389;
	assign origtmp1824 = in[1219] ^ origtmp1737;
	assign origtmp1820 = origtmp1805 ^ in[427];
	assign origtmp476 = in[738] ^ origtmp475;
	assign out[430] = 1'b0 & 1'b0;
	assign origtmp1417 = origtmp1910 ^ origtmp1672;
	assign origtmp220 = origtmp218;
	assign origtmp638 = 1'b1 | 1'b1;
	assign origtmp2222 = in[1132] & origtmp1452;
	assign origtmp1476 = in[177] | in[760];
	assign origtmp821 = ~origtmp820;
	assign origtmp2103 = origtmp1998 & in[921];
	assign out[484] = ~in[564];
	assign origtmp459 = origtmp460 ^ origtmp462;
	assign origtmp197 = origtmp199 ^ origtmp198;
	assign origtmp1075 = 1'b1 & in[957];
	assign origtmp1662 = in[259] & in[184];
	assign origtmp595 = in[1236] & origtmp596;
	assign origtmp1809 = origtmp2047 | in[483];
	assign out[213] = origtmp525 ^ origtmp527;
	assign origtmp324 = origtmp325 ^ origtmp325;
	assign origtmp1951 = origtmp1480 ^ origtmp1361;
	assign out[109] = in[458] ^ in[458];
	assign origtmp1440 = in[914] ^ origtmp1696;
	assign origtmp105 = origtmp106 & origtmp107;
	assign origtmp298 = in[737] | 1'b1;
	assign origtmp115 = 1'b1;
	assign origtmp1735 = in[917] | origtmp1886;
	assign origtmp1295 = origtmp1748 | in[95];
	assign origtmp1464 = in[178] & in[871];
	assign origtmp2026 = in[1396] ^ origtmp1340;
	assign out[389] = origtmp962 | origtmp963;
	assign out[361] = origtmp898 ^ origtmp897;
	assign origtmp282 = 1'b0 | 1'b1;
	assign out[23] = origtmp60 ^ in[330];
	assign origtmp233 = origtmp232 | 1'b1;
	assign origtmp2033 = in[470] | in[127];
	assign origtmp318 = ~origtmp319;
	assign origtmp904 = 1'b0;
	assign out[340] = 1'b0 ^ origtmp849;
	assign origtmp1995 = origtmp1256 ^ in[773];
	assign origtmp1801 = in[790] | in[1428];
	assign origtmp2054 = origtmp1645 & in[89];
	assign origtmp1729 = origtmp2132 ^ in[234];
	assign origtmp1155 = origtmp1152 ^ origtmp1152;
	assign origtmp1364 = in[858] | in[323];
	assign origtmp77 = ~1'b1;
	assign origtmp669 = in[1100];
	assign origtmp16 = in[823] ^ 1'b1;
	assign origtmp307 = 1'b1 | 1'b0;
	assign origtmp242 = 1'b0 ^ origtmp244;
	assign origtmp142 = in[289] ^ 1'b0;
	assign origtmp1387 = in[1145] ^ in[1019];
	assign origtmp697 = in[1157] & in[976];
	assign origtmp896 = origtmp895 & origtmp894;
	assign origtmp455 = 1'b0 & 1'b0;
	assign origtmp6 = in[1486] | origtmp7;
	assign out[38] = origtmp99 ^ 1'b1;
	assign origtmp1175 = origtmp1176 | origtmp1176;
	assign origtmp325 = 1'b0 & in[1117];
	assign origtmp432 = in[539];
	assign origtmp2143 = origtmp1367 & in[1381];
	assign origtmp1675 = in[191] | in[4];
	assign origtmp491 = origtmp493 | 1'b0;
	assign out[171] = origtmp428 ^ origtmp431;
	assign origtmp1120 = origtmp1122 & 1'b1;
	assign origtmp398 = origtmp399;
	assign origtmp1247 = in[394] ^ in[546];
	assign origtmp1133 = 1'b0 ^ 1'b0;
	assign origtmp840 = origtmp841 ^ 1'b1;
	assign origtmp2252 = origtmp1442 | origtmp1445;
	assign origtmp1358 = origtmp1756 & origtmp1308;
	assign origtmp2016 = in[1148] ^ in[302];
	assign origtmp1782 = origtmp2052 | origtmp1883;
	assign origtmp32 = origtmp36 | 1'b1;
	assign origtmp938 = 1'b1 | 1'b1;
	assign origtmp1778 = origtmp1648 ^ origtmp1715;
	assign origtmp893 = origtmp892 | 1'b0;
	assign origtmp2158 = origtmp2161 ^ in[15];
	assign origtmp37 = 1'b0 | 1'b1;
	assign origtmp296 = in[1403] ^ in[973];
	assign out[12] = in[1379] | in[1366];
	assign origtmp279 = 1'b1 & 1'b1;
	assign origtmp63 = 1'b1 & in[1334];
	assign origtmp1486 = in[54] & origtmp2008;
	assign origtmp1621 = in[135] ^ in[176];
	assign origtmp2246 = origtmp1320 | origtmp2163;
	assign origtmp766 = in[151] | 1'b1;
	assign origtmp1560 = origtmp1996 & origtmp2101;
	assign out[245] = origtmp607 & origtmp608;
	assign origtmp423 = origtmp426 | in[35];
	assign origtmp1178 = origtmp1179 | 1'b1;
	assign out[181] = origtmp448;
	assign origtmp1083 = 1'b0;
	assign origtmp1550 = origtmp2137 ^ origtmp2116;
	assign origtmp1581 = in[253] ^ origtmp1920;
	assign origtmp1221 = ~in[240];
	assign origtmp489 = 1'b1 & origtmp488;
	assign origtmp2125 = in[561] | origtmp1517;
	assign origtmp946 = origtmp943 ^ origtmp943;
	assign origtmp1452 = origtmp1323 | in[482];
	assign origtmp368 = in[828] & origtmp369;
	assign origtmp1212 = origtmp1210 & origtmp1210;
	assign origtmp990 = origtmp988 & 1'b1;
	assign origtmp1641 = origtmp2100 & origtmp1786;
	assign origtmp574 = ~1'b1;
	assign origtmp393 = in[583] & origtmp391;
	assign origtmp85 = origtmp83 | in[123];
	assign origtmp76 = 1'b1 & in[1364];
	assign origtmp1274 = in[612] | in[377];
	assign out[413] = origtmp1013 | in[72];
	assign origtmp1034 = in[1202] & in[1202];
	assign origtmp961 = origtmp960 ^ in[230];
	assign out[81] = origtmp197;
	assign origtmp721 = origtmp720 ^ origtmp719;
	assign origtmp1007 = in[1363] | 1'b1;
	assign origtmp1148 = 1'b0 & origtmp1150;
	assign out[82] = origtmp205 ^ origtmp202;
	assign origtmp940 = in[551];
	assign origtmp1135 = in[1104] | origtmp1137;
	assign origtmp1507 = in[214] & origtmp1684;
	assign origtmp1882 = origtmp1300 ^ origtmp1390;
	assign origtmp1619 = in[1170] & origtmp1721;
	assign out[463] = in[554] ^ origtmp1163;
	assign origtmp1112 = ~1'b0;
	assign origtmp88 = origtmp89 | 1'b1;
	assign out[390] = in[874] & origtmp964;
	assign origtmp1925 = in[890] ^ origtmp1771;
	assign origtmp531 = in[203] & in[339];
	assign origtmp2124 = in[371] | in[1301];
	assign out[204] = in[480] ^ origtmp514;
	assign origtmp933 = 1'b0 ^ 1'b0;
	assign origtmp1939 = in[1445] | origtmp1577;
	assign origtmp1947 = in[1355] | in[1193];
	assign origtmp253 = in[1133] & in[1099];
	assign origtmp249 = origtmp250 | origtmp248;
	assign origtmp1139 = in[156];
	assign origtmp1480 = origtmp1804 | origtmp1671;
	assign origtmp2005 = in[722] ^ origtmp1609;
	assign origtmp885 = origtmp886 | origtmp887;
	assign out[176] = ~1'b0;
	assign origtmp1512 = origtmp1699 | origtmp1936;
	assign origtmp1692 = origtmp2168 ^ origtmp1911;
	assign origtmp607 = 1'b1 | origtmp609;
	assign origtmp1726 = in[1370] & in[42];
	assign out[448] = origtmp1114 & origtmp1113;
	assign origtmp1261 = origtmp1923 & origtmp2057;
	assign origtmp1865 = in[1015] | in[466];
	assign origtmp1914 = in[395] & in[656];
	assign origtmp355 = 1'b1 & origtmp356;
	assign out[193] = 1'b0 ^ origtmp484;
	assign origtmp276 = origtmp274 | 1'b1;
	assign origtmp826 = origtmp824;
	assign out[375] = origtmp924;
	assign origtmp1698 = in[223] ^ origtmp1476;
	assign origtmp322 = origtmp323 | 1'b0;
	assign origtmp758 = 1'b0;
	assign origtmp2112 = in[287] ^ origtmp1499;
	assign origtmp1081 = origtmp1082 & origtmp1083;
	assign origtmp500 = 1'b1 ^ origtmp503;
	assign origtmp217 = 1'b1 ^ 1'b1;
	assign out[488] = 1'b1 & origtmp1219;
	assign origtmp716 = 1'b1 ^ in[562];
	assign out[462] = 1'b0 & origtmp1160;
	assign origtmp1058 = origtmp1059 & 1'b0;
	assign origtmp625 = ~origtmp626;
	assign origtmp1708 = in[866] | in[1471];
	assign origtmp310 = ~1'b0;
	assign origtmp1904 = in[1433] | origtmp1675;
	assign origtmp1724 = in[469] & in[573];
	assign origtmp1658 = in[278] & origtmp2050;
	assign origtmp1797 = in[1048] & in[322];
	assign out[400] = origtmp992 & origtmp993;
	assign origtmp1953 = in[615] | in[1211];
	assign origtmp1211 = in[1400] | in[649];
	assign out[235] = 1'b1 & 1'b0;
	assign origtmp315 = 1'b0 | in[98];
	assign origtmp2097 = in[657] ^ in[801];
	assign origtmp1269 = origtmp1631 | in[1109];
	assign origtmp1450 = in[450] & in[755];
	assign origtmp2071 = origtmp2025 ^ origtmp2236;
	assign origtmp1847 = in[616] | origtmp1809;
	assign origtmp190 = in[439] ^ 1'b1;
	assign origtmp709 = ~1'b0;
	assign origtmp192 = 1'b0 | 1'b1;
	assign origtmp441 = ~in[560];
	assign out[215] = origtmp532 ^ 1'b1;
	assign out[416] = origtmp1025 ^ origtmp1023;
	assign origtmp236 = 1'b1 ^ in[1074];
	assign origtmp2023 = origtmp1742 ^ origtmp1369;
	assign out[297] = 1'b0;
	assign origtmp229 = ~in[676];
	assign origtmp927 = origtmp925 ^ origtmp926;
	assign origtmp208 = origtmp211 & 1'b0;
	assign origtmp1165 = origtmp1164 & origtmp1164;
	assign out[248] = origtmp619 ^ origtmp617;
	assign origtmp314 = ~origtmp315;
	assign origtmp685 = 1'b0;
	assign origtmp2086 = origtmp1719 & origtmp2070;
	assign origtmp1288 = origtmp1572 & in[75];
	assign origtmp258 = origtmp260 | origtmp259;
	assign origtmp732 = origtmp734 | in[767];
	assign out[490] = origtmp1224 ^ origtmp1224;
	assign origtmp1369 = in[307] & in[1221];
	assign origtmp1751 = in[1372] & in[231];
	assign origtmp1224 = 1'b1;
	assign origtmp1381 = in[499] | in[527];
	assign origtmp171 = 1'b0 & 1'b0;
	assign origtmp1543 = in[1116] ^ origtmp2152;
	assign origtmp839 = in[702] & in[1254];
	assign origtmp1558 = origtmp1693 & origtmp2005;
	assign origtmp516 = in[894] | in[1255];
	assign origtmp1572 = origtmp1348 | in[1481];
	assign out[330] = in[432] | in[341];
	assign origtmp1671 = origtmp1857 | origtmp1302;
	assign origtmp1601 = origtmp1521 ^ origtmp2188;
	assign origtmp930 = origtmp931 & in[981];
	assign out[454] = origtmp1134 & origtmp1136;
	assign origtmp1094 = origtmp1095 ^ 1'b1;
	assign out[67] = origtmp171 | origtmp172;
	assign origtmp269 = in[569] & 1'b1;
	assign origtmp1065 = origtmp1066 | origtmp1066;
	assign origtmp573 = ~origtmp574;
	assign origtmp1305 = in[768] | in[171];
	assign origtmp1304 = origtmp2016 & in[1144];
	assign origtmp1715 = origtmp2233 & origtmp1852;
	assign origtmp440 = in[74] ^ in[74];
	assign origtmp2179 = in[1055] ^ in[1304];
	assign out[28] = origtmp76 ^ in[1364];
	assign out[122] = 1'b0 ^ origtmp303;
	assign origtmp1967 = in[1238] | in[869];
	assign origtmp1689 = in[766] ^ in[948];
	assign origtmp684 = origtmp685 & origtmp686;
	assign out[44] = in[1077] & in[807];
	assign origtmp1762 = in[912] & in[928];
	assign origtmp2089 = in[375] & in[362];
	assign out[11] = origtmp27 ^ 1'b1;
	assign origtmp486 = 1'b1;
	assign origtmp1978 = origtmp1613 & in[1469];
	assign origtmp434 = origtmp436 | in[539];
	assign out[422] = origtmp1043 | origtmp1044;
	assign out[177] = origtmp442 & origtmp441;
	assign out[76] = origtmp189 & origtmp189;
	assign out[75] = in[1453] | origtmp188;
	assign origtmp1293 = in[225] | origtmp1363;
	assign origtmp723 = origtmp722 & in[208];
	assign origtmp1607 = origtmp1764 | origtmp1514;
	assign origtmp1123 = 1'b0 | in[273];
	assign origtmp57 = ~1'b0;
	assign origtmp1190 = origtmp1188 & origtmp1188;
	assign out[56] = origtmp138 ^ origtmp138;
	assign origtmp1203 = 1'b1 | 1'b0;
	assign out[161] = origtmp403 | origtmp403;
	assign origtmp901 = in[1299] | 1'b1;
	assign origtmp764 = in[784] ^ in[151];
	assign origtmp2235 = origtmp1578 | origtmp1922;
	assign origtmp1763 = origtmp2201 & in[103];
	assign origtmp155 = 1'b1 ^ origtmp154;
	assign origtmp751 = 1'b0 ^ 1'b0;
	assign origtmp2061 = origtmp1677 | origtmp1723;
	assign origtmp2075 = origtmp1826 ^ origtmp1979;
	assign origtmp2148 = origtmp1241 & origtmp2243;
	assign origtmp701 = origtmp702 & 1'b1;
	assign origtmp1016 = origtmp1015 ^ origtmp1015;
	assign origtmp1402 = in[1013] | in[970];
	assign origtmp264 = 1'b0 | origtmp262;
	assign out[73] = origtmp182 | 1'b0;
	assign origtmp1053 = 1'b1;
	assign origtmp1871 = in[591] | in[413];
	assign origtmp9 = in[383] ^ in[1474];
	assign origtmp1037 = origtmp1038 | origtmp1036;
	assign out[256] = origtmp634 ^ origtmp636;
	assign out[126] = in[365];
	assign out[211] = in[1172] | origtmp520;
	assign origtmp1275 = in[1095] ^ in[1464];
	assign origtmp1185 = origtmp1184 ^ 1'b0;
	assign origtmp1875 = origtmp2020 ^ origtmp1966;
	assign origtmp952 = 1'b1 | origtmp954;
	assign origtmp1096 = in[524] ^ origtmp1092;
	assign origtmp91 = origtmp93 ^ 1'b0;
	assign origtmp1659 = in[34] | in[281];
	assign origtmp2133 = origtmp1388 ^ origtmp2121;
	assign out[326] = 1'b0 | origtmp809;
	assign out[358] = origtmp893 ^ 1'b0;
	assign origtmp1383 = in[1386] | origtmp2185;
	assign origtmp2046 = in[959] & origtmp1977;
	assign origtmp796 = origtmp797 ^ origtmp797;
	assign out[364] = origtmp902 ^ origtmp903;
	assign origtmp1365 = origtmp1279 & origtmp1991;
	assign origtmp1035 = 1'b1 | 1'b0;
	assign out[440] = origtmp1089 ^ origtmp1090;
	assign origtmp1717 = origtmp2072 | origtmp1317;
	assign out[486] = in[927] & in[1204];
	assign origtmp1712 = in[1398] | origtmp1788;
	assign origtmp1599 = origtmp2107 | origtmp2098;
	assign origtmp2245 = in[1297] & origtmp1623;
	assign origtmp2118 = origtmp1415 | origtmp1346;
	assign origtmp802 = origtmp804;
	assign out[266] = origtmp662 ^ origtmp664;
	assign out[229] = origtmp576 & origtmp575;
	assign origtmp887 = origtmp888;
	assign out[294] = origtmp744 ^ in[944];
	assign origtmp400 = in[772] | 1'b0;
	assign origtmp2177 = in[213] ^ origtmp1259;
	assign origtmp1020 = 1'b1 ^ origtmp1019;
	assign origtmp1876 = in[1275] & origtmp1561;
	assign origtmp1259 = in[441] ^ in[533];
	assign origtmp1367 = in[167] | in[876];
	assign origtmp2130 = in[1483] & in[929];
	assign origtmp2098 = origtmp2166 | origtmp1385;
	assign origtmp779 = ~origtmp780;
	assign origtmp1197 = in[660];
	assign out[226] = origtmp568 & 1'b1;
	assign origtmp56 = 1'b0 ^ 1'b0;
	assign origtmp1268 = origtmp1896 & origtmp1959;
	assign out[404] = 1'b0 & origtmp998;
	assign origtmp823 = in[210] | origtmp821;
	assign origtmp829 = in[833] & 1'b0;
	assign origtmp1990 = origtmp1536 & origtmp1258;
	assign out[385] = origtmp947 | origtmp948;
	assign origtmp367 = origtmp368 ^ in[1387];
	assign origtmp1057 = origtmp1059 & origtmp1058;
	assign origtmp449 = origtmp450 ^ 1'b1;
	assign out[397] = 1'b0 & origtmp984;
	assign origtmp1589 = origtmp1639 & in[555];
	assign origtmp1378 = origtmp2028 | origtmp2089;
	assign origtmp1285 = in[611] | origtmp1359;
	assign out[387] = 1'b1 & 1'b1;
	assign origtmp2110 = origtmp1269 | origtmp1697;
	assign origtmp1503 = in[968] | in[1418];
	assign out[436] = origtmp1081 & origtmp1084;
	assign origtmp2031 = origtmp1787 | in[540];
	assign origtmp1626 = in[1472] ^ origtmp1685;
	assign origtmp82 = in[123];
	assign origtmp1029 = 1'b0 & origtmp1027;
	assign out[63] = origtmp158 | in[872];
	assign origtmp193 = 1'b0;
	assign origtmp1804 = in[559] | origtmp1855;
	assign origtmp1116 = 1'b1 ^ in[266];
	assign origtmp730 = 1'b1;
	assign origtmp724 = origtmp722 ^ origtmp723;
	assign origtmp875 = 1'b1 ^ origtmp874;
	assign origtmp555 = origtmp554 & in[479];
	assign origtmp727 = origtmp728 | in[274];
	assign origtmp1436 = in[1286] | in[750];
	assign out[234] = in[10] | in[201];
	assign origtmp445 = origtmp444 & origtmp444;
	assign origtmp1841 = origtmp2190 & in[1014];
	assign origtmp1817 = origtmp1836 | in[854];
	assign origtmp178 = origtmp179 ^ in[558];
	assign origtmp1283 = origtmp1651 ^ in[1022];
	assign origtmp327 = origtmp326;
	assign out[192] = origtmp479 & origtmp480;
	assign origtmp540 = 1'b0 & 1'b0;
	assign out[218] = origtmp542 | origtmp544;
	assign origtmp1177 = 1'b0 & in[600];
	assign origtmp399 = 1'b1 | in[772];
	assign origtmp133 = in[1032] ^ 1'b1;
	assign origtmp477 = 1'b0 & 1'b0;
	assign out[6] = in[1196] | 1'b1;
	assign origtmp1055 = origtmp1056 & origtmp1054;
	assign origtmp1439 = origtmp2235 ^ origtmp1660;
	assign origtmp655 = 1'b0;
	assign origtmp1401 = origtmp1860 & origtmp1867;
	assign origtmp639 = ~1'b0;
	assign origtmp813 = origtmp812 ^ origtmp811;
	assign origtmp1086 = in[1178] ^ 1'b0;
	assign origtmp1897 = origtmp1554 & origtmp1683;
	assign origtmp747 = origtmp750 & origtmp750;
	assign origtmp1374 = in[1112] & in[528];
	assign origtmp1553 = in[1457] | origtmp2051;
	assign origtmp1654 = in[724] | in[1371];
	assign origtmp2211 = origtmp1610 | in[1312];
	assign origtmp811 = in[1332] & origtmp810;
	assign out[43] = origtmp112 ^ origtmp111;
	assign origtmp1509 = origtmp1291 & origtmp2212;
	assign origtmp1208 = origtmp1204 ^ origtmp1205;
	assign origtmp994 = in[1106] & in[53];
	assign origtmp333 = 1'b1 ^ 1'b1;
	assign out[270] = origtmp675 ^ 1'b1;
	assign origtmp1117 = origtmp1118 & in[541];
	assign origtmp680 = 1'b0 & 1'b0;
	assign origtmp391 = in[709];
	assign out[111] = origtmp279 | origtmp280;
	assign origtmp1860 = in[608] & in[908];
	assign origtmp1006 = origtmp1004 & 1'b0;
	assign out[481] = ~1'b1;
	assign out[362] = origtmp900 & 1'b1;
	assign out[338] = origtmp843 & origtmp842;
	assign origtmp776 = origtmp775 & 1'b0;
	assign origtmp683 = 1'b1 & origtmp684;
	assign origtmp1975 = in[279] ^ in[1136];
	assign origtmp48 = origtmp51 ^ in[905];
	assign origtmp1518 = origtmp1733 ^ origtmp2162;
	assign origtmp64 = ~1'b0;
	assign origtmp1219 = 1'b1 ^ origtmp1223;
	assign origtmp1937 = in[498] ^ origtmp1665;
	assign origtmp188 = ~origtmp187;
	assign origtmp1551 = in[212] | origtmp1380;
	assign origtmp1229 = in[79] | 1'b1;
	assign origtmp98 = 1'b1 | origtmp97;
	assign origtmp1810 = origtmp1806 | in[282];
	assign out[443] = in[1258] & origtmp1098;
	assign out[344] = ~in[491];
	assign origtmp1677 = origtmp1573 | origtmp2157;
	assign origtmp1171 = 1'b1 & in[1246];
	assign origtmp664 = origtmp665 | origtmp665;
	assign origtmp2147 = origtmp1565 & origtmp1624;
	assign origtmp2050 = in[875] ^ origtmp1253;
	assign origtmp1575 = in[68] ^ in[1186];
	assign out[367] = 1'b0 & origtmp906;
	assign origtmp1792 = in[563] ^ origtmp1513;
	assign origtmp593 = 1'b0;
	assign origtmp1709 = in[685] & in[580];
	assign origtmp216 = 1'b1 ^ origtmp213;
	assign origtmp1757 = in[961] & in[1368];
	assign origtmp749 = 1'b1 ^ 1'b1;
	assign origtmp54 = origtmp57 | 1'b1;
	assign origtmp438 = ~1'b1;
	assign origtmp1172 = ~origtmp1171;
	assign out[119] = 1'b0 & origtmp296;
	assign origtmp113 = in[701] | in[870];
	assign origtmp622 = 1'b1 & 1'b1;
	assign origtmp1428 = in[1184] | in[325];
	assign origtmp1750 = in[506] & origtmp1746;
	assign origtmp451 = 1'b0 & 1'b0;
	assign origtmp611 = in[57] & origtmp610;
	assign origtmp1613 = origtmp1426 & in[308];
	assign origtmp1121 = origtmp1124 & in[273];
	assign origtmp273 = origtmp275 ^ in[387];
	assign out[112] = origtmp282 ^ origtmp283;
	assign origtmp2020 = in[180] & in[101];
	assign out[72] = origtmp178 & in[1426];
	assign origtmp2173 = in[1149] & origtmp1628;
	assign origtmp1144 = in[328] ^ origtmp1142;
	assign out[42] = origtmp108 ^ origtmp109;
	assign origtmp2228 = origtmp2088 ^ origtmp1409;
	assign origtmp1857 = origtmp2250 | origtmp1644;
	assign origtmp2105 = in[845] ^ origtmp2248;
	assign origtmp260 = in[1188] & in[1188];
	assign origtmp1610 = origtmp1596 & origtmp1475;
	assign origtmp388 = origtmp387 | origtmp387;
	assign origtmp244 = 1'b0;
	assign origtmp1772 = origtmp1364 | origtmp1755;
	assign origtmp587 = 1'b1 | in[1272];
	assign origtmp1540 = in[60] | origtmp1728;
	assign origtmp1189 = 1'b0 | origtmp1190;
	assign origtmp817 = origtmp815 | in[748];
	assign origtmp1011 = 1'b0;
	assign origtmp1625 = origtmp1293 & origtmp2175;
	assign origtmp621 = in[1115] & 1'b0;
	assign origtmp1948 = in[646] & origtmp1667;
	assign origtmp1513 = in[1182] & in[118];
	assign origtmp1316 = origtmp1266 | origtmp1263;
	assign origtmp895 = in[1447] | in[804];
	assign origtmp842 = 1'b1;
	assign origtmp1595 = origtmp1868 ^ in[250];
	assign origtmp1508 = origtmp2026 | origtmp2031;
	assign origtmp419 = ~origtmp421;
	assign origtmp2115 = in[1348] ^ origtmp1814;
	assign origtmp1386 = origtmp1650 & origtmp1952;
	assign origtmp2206 = in[476] ^ origtmp1487;
	assign out[284] = origtmp721 ^ origtmp718;
	assign origtmp1469 = in[128] ^ origtmp1726;
	assign origtmp2214 = in[1129] ^ origtmp2041;
	assign origtmp1908 = in[1322] ^ in[64];
	assign origtmp2242 = origtmp1358 ^ origtmp2073;
	assign out[223] = origtmp558 & origtmp561;
	assign origtmp302 = 1'b1 ^ 1'b1;
	assign origtmp39 = origtmp40 | 1'b0;
	assign origtmp1915 = in[1284] ^ in[111];
	assign out[377] = origtmp930 & in[33];
	assign out[483] = origtmp1213 ^ origtmp1212;
	assign origtmp1821 = origtmp1280 | origtmp2075;
	assign origtmp1167 = 1'b1 & 1'b1;
	assign origtmp2239 = in[142] & in[919];
	assign origtmp174 = origtmp176 & 1'b0;
	assign out[499] = origtmp1663 & origtmp1391;
	assign origtmp909 = in[316] | origtmp908;
	assign origtmp2079 = origtmp1336 ^ origtmp1337;
	assign origtmp70 = 1'b1;
	assign origtmp799 = 1'b0 & origtmp798;
	assign origtmp917 = origtmp916 ^ in[168];
	assign origtmp910 = origtmp912 | in[1264];
	assign out[359] = 1'b0 ^ origtmp896;
	assign origtmp1141 = origtmp1140 & origtmp1139;
	assign out[325] = 1'b1 | origtmp808;
	assign out[207] = origtmp515 | 1'b0;
	assign out[143] = 1'b1 | 1'b0;
	assign origtmp40 = origtmp42 ^ 1'b1;
	assign origtmp1919 = origtmp1443 | origtmp2154;
	assign origtmp586 = 1'b1 ^ 1'b1;
	assign out[347] = in[926] & in[298];
	assign out[27] = in[1295] & origtmp75;
	assign origtmp1388 = origtmp1347 & in[1085];
	assign origtmp1668 = origtmp1942 | in[512];
	assign origtmp756 = in[1171] & in[1171];
	assign origtmp362 = ~1'b0;
	assign origtmp26 = origtmp22 | 1'b1;
	assign origtmp319 = 1'b0 & in[1268];
	assign origtmp297 = in[1417];
	assign origtmp1534 = in[689] & origtmp1276;
	assign origtmp1337 = in[1029] | origtmp2043;
	assign out[285] = ~in[534];
	assign out[103] = origtmp258 ^ origtmp257;
	assign origtmp337 = in[1335] ^ origtmp339;
	assign origtmp2091 = in[638] & in[14];
	assign origtmp1670 = in[831] & in[1153];
	assign origtmp1100 = ~1'b1;
	assign origtmp374 = in[48] ^ in[48];
	assign origtmp1420 = in[449] & in[190];
	assign origtmp600 = 1'b1 ^ origtmp601;
	assign origtmp376 = in[1002] | origtmp372;
	assign origtmp2167 = in[428] ^ in[1228];
	assign origtmp871 = origtmp873;
	assign origtmp163 = ~in[320];
	assign origtmp414 = origtmp417 & origtmp418;
	assign out[49] = origtmp121 ^ origtmp119;
	assign origtmp185 = 1'b0 | in[20];
	assign origtmp1416 = in[855] & in[200];
	assign origtmp1781 = in[1247] ^ origtmp1474;
	assign origtmp184 = 1'b1 & origtmp183;
	assign origtmp379 = origtmp377 & origtmp377;
	assign out[496] = in[136] | origtmp1234;
	assign origtmp2087 = origtmp1617 | origtmp1508;
	assign origtmp4 = 1'b0 ^ 1'b1;
	assign origtmp1800 = origtmp1619 ^ origtmp1612;
	assign out[319] = origtmp793 ^ origtmp794;
	assign origtmp1340 = in[1189] & in[1165];
	assign out[100] = 1'b0 | origtmp251;
	assign origtmp493 = ~1'b1;
	assign origtmp618 = in[131] | 1'b0;
	assign origtmp410 = origtmp412 & origtmp411;
	assign origtmp1731 = origtmp2007 ^ in[566];
	assign origtmp2047 = in[793] & in[667];
	assign out[475] = origtmp1193 & origtmp1194;
	assign out[163] = 1'b0 | origtmp409;
	assign out[292] = 1'b1 | 1'b1;
	assign out[101] = origtmp253 & in[1133];
	assign out[282] = origtmp709 | origtmp712;
	assign out[357] = origtmp890 & origtmp891;
	assign origtmp65 = in[952] ^ 1'b1;
	assign out[276] = origtmp693 & origtmp695;
	assign origtmp1591 = origtmp1257 ^ origtmp1845;
	assign out[107] = origtmp272 | origtmp270;
	assign origtmp469 = in[644] ^ 1'b0;
	assign origtmp2178 = origtmp2173 | origtmp1939;
	assign origtmp1886 = in[710] | in[899];
	assign origtmp14 = origtmp16 ^ 1'b1;
	assign out[371] = origtmp913 ^ origtmp914;
	assign out[190] = origtmp474 ^ 1'b0;
	assign origtmp1000 = 1'b1;
	assign origtmp1548 = origtmp1642 ^ origtmp1717;
	assign out[59] = 1'b1 & origtmp145;
	assign origtmp771 = origtmp769 | origtmp769;
	assign origtmp1251 = origtmp1355 | origtmp1261;
	assign out[498] = origtmp1238 ^ origtmp1239;
	assign origtmp1366 = in[792] | in[1444];
	assign origtmp2218 = origtmp2093 | in[226];
	assign origtmp921 = 1'b0 ^ origtmp923;
	assign origtmp1406 = origtmp1766 ^ in[619];
	assign origtmp792 = 1'b1;
	assign origtmp1142 = 1'b0 & in[328];
	assign origtmp2095 = in[1147] | origtmp2125;
	assign origtmp1687 = in[1408] | in[1475];
	assign origtmp1501 = origtmp1547 | origtmp1915;
	assign origtmp2055 = origtmp2148 & origtmp2221;
	assign origtmp918 = 1'b0 | origtmp919;
	assign origtmp1505 = in[244] | in[398];
	assign origtmp168 = origtmp170 & origtmp170;
	assign out[212] = 1'b0 & origtmp523;
	assign origtmp1565 = in[607] ^ origtmp1366;
	assign origtmp1336 = in[1028] | origtmp2109;
	assign origtmp1853 = in[1231] | origtmp2063;
	assign origtmp1325 = in[1159] & in[485];
	assign origtmp484 = origtmp483 | origtmp482;
	assign origtmp743 = in[235] | 1'b0;
	assign origtmp905 = ~in[29];
	assign origtmp149 = 1'b1;
	assign origtmp1355 = origtmp1669 | origtmp1661;
	assign out[97] = origtmp247 & origtmp246;
	assign origtmp903 = 1'b1;
	assign origtmp2114 = in[730] & origtmp1891;
	assign origtmp331 = ~origtmp330;
	assign origtmp1828 = origtmp1777 ^ origtmp1918;
	assign origtmp448 = 1'b0 ^ in[115];
	assign origtmp415 = in[255] & in[255];
	assign origtmp1685 = in[575] ^ origtmp1908;
	assign origtmp104 = 1'b1 & in[933];
	assign origtmp636 = ~in[130];
	assign out[167] = in[1127] | 1'b1;
	assign out[383] = 1'b0 ^ origtmp942;
	assign origtmp34 = ~1'b1;
	assign origtmp499 = in[549] ^ 1'b0;
	assign out[467] = origtmp1169 ^ origtmp1173;
	assign origtmp79 = origtmp81;
	assign origtmp1079 = in[414];
	assign out[128] = origtmp322 | origtmp321;
	assign origtmp1979 = origtmp2082 & origtmp1901;
	assign origtmp62 = origtmp64;
	assign out[250] = origtmp624 | origtmp622;
	assign origtmp1696 = in[915] ^ in[988];
	assign origtmp582 = in[1276] ^ in[775];
	assign origtmp128 = 1'b1 | in[1338];
	assign origtmp892 = ~1'b0;
	assign origtmp1270 = origtmp1793 ^ origtmp2147;
	assign origtmp950 = 1'b1 ^ 1'b1;
	assign origtmp1110 = origtmp1111 ^ origtmp1111;
	assign origtmp1635 = origtmp2079 | in[542];
	assign origtmp1639 = in[59] & in[743];
	assign out[352] = in[486] & origtmp877;
	assign origtmp1905 = origtmp1821 & origtmp2102;
	assign origtmp2080 = in[27] ^ in[437];
	assign origtmp715 = ~origtmp716;
	assign out[186] = origtmp459 | origtmp461;
	assign origtmp535 = 1'b0;
	assign origtmp2186 = in[454] | origtmp2209;
	assign origtmp1665 = origtmp1797 ^ in[980];
	assign origtmp2077 = in[447] & in[1411];
	assign origtmp1382 = origtmp1314 ^ origtmp2189;
	assign origtmp1765 = origtmp1992 ^ origtmp1534;
	assign origtmp1179 = origtmp1180 ^ origtmp1181;
	assign origtmp1384 = in[879] | origtmp1862;
	assign origtmp1004 = 1'b1;
	assign origtmp882 = origtmp880 ^ in[1010];
	assign out[335] = origtmp837 | 1'b1;
	assign origtmp1363 = in[66] | origtmp1535;
	assign origtmp1243 = origtmp1462 | origtmp1828;
	assign origtmp2199 = in[76] & in[622];
	assign origtmp2014 = in[349] ^ in[1307];
	assign out[144] = origtmp357 & origtmp355;
	assign origtmp1485 = in[452] & in[28];
	assign origtmp1785 = in[489] | in[759];
	assign origtmp1348 = in[25] ^ origtmp1360;
	assign origtmp967 = ~1'b1;
	assign origtmp1026 = origtmp1028 & origtmp1029;
	assign origtmp596 = in[1236];
	assign out[180] = origtmp447 | origtmp446;
	assign origtmp757 = origtmp756 & origtmp755;
	assign origtmp212 = 1'b1 & 1'b1;
	assign origtmp851 = 1'b1 & origtmp852;
	assign origtmp1693 = in[1083] ^ in[824];
	assign origtmp2123 = origtmp2015 ^ origtmp2172;
	assign origtmp929 = origtmp928 & origtmp927;
	assign origtmp1922 = origtmp1601 | origtmp1951;
	assign out[196] = 1'b0 | origtmp492;
	assign origtmp1917 = in[1195] & origtmp1588;
	assign origtmp2141 = in[248] | in[1434];
	assign origtmp1956 = in[1288] & in[1282];
	assign origtmp238 = origtmp237 | origtmp239;
	assign origtmp1113 = origtmp1112 ^ 1'b1;
	assign origtmp633 = in[503] | in[1007];
	assign origtmp139 = ~in[1018];
	assign out[24] = origtmp62 | origtmp61;
	assign origtmp151 = 1'b1;
	assign origtmp603 = origtmp600 ^ origtmp602;
	assign origtmp162 = 1'b1;
	assign origtmp578 = 1'b1;
	assign origtmp934 = origtmp933 | origtmp935;
	assign origtmp74 = ~1'b1;
	assign origtmp1279 = origtmp2076 | origtmp2192;
	assign out[402] = origtmp996 ^ origtmp995;
	assign out[314] = in[310] & origtmp787;
	assign origtmp705 = 1'b0 | origtmp704;
	assign origtmp1054 = 1'b1 ^ origtmp1053;
	assign origtmp1921 = in[645] & in[813];
	assign origtmp1360 = origtmp2226 & in[693];
	assign origtmp713 = 1'b1 | in[846];
	assign out[87] = origtmp220 & origtmp219;
	assign out[52] = origtmp130 & origtmp129;
	assign origtmp1095 = origtmp1093 ^ in[524];
	assign origtmp590 = origtmp592 ^ origtmp593;
	assign out[343] = in[651] ^ in[825];
	assign out[355] = origtmp885 | origtmp885;
	assign origtmp602 = 1'b1 ^ origtmp604;
	assign origtmp1739 = origtmp1463 | origtmp1576;
	assign origtmp1652 = origtmp1512 & origtmp2145;
	assign origtmp289 = 1'b0 | 1'b0;
	assign origtmp294 = 1'b1;
	assign origtmp514 = 1'b0 | in[1240];
	assign out[293] = origtmp742 | origtmp741;
	assign origtmp1196 = origtmp1198 | 1'b1;
	assign origtmp173 = origtmp176;
	assign origtmp1720 = in[1056] | in[206];
	assign origtmp259 = in[1188] & in[670];
	assign origtmp644 = origtmp645 & 1'b1;
	assign origtmp682 = in[207] | 1'b0;
	assign origtmp1971 = origtmp1362 ^ origtmp1498;
	assign origtmp473 = origtmp469 ^ 1'b0;
	assign origtmp1633 = in[456] & origtmp1708;
	assign origtmp442 = in[97];
	assign origtmp1435 = in[1050] | in[553];
	assign out[480] = origtmp1207 & origtmp1208;
	assign out[150] = origtmp373 ^ origtmp375;
	assign origtmp2 = origtmp3 | 1'b1;
	assign origtmp854 = 1'b0 & 1'b1;
	assign out[10] = origtmp23 ^ origtmp24;
	assign origtmp2094 = in[826] | in[637];
	assign origtmp116 = ~origtmp117;
	assign out[445] = origtmp1107 ^ origtmp1105;
	assign origtmp100 = in[504] | in[504];
	assign out[19] = origtmp48 ^ origtmp49;
	assign origtmp153 = 1'b0;
	assign out[160] = origtmp401 | 1'b1;
	assign origtmp1858 = origtmp1435 ^ origtmp1854;
	assign origtmp2074 = origtmp1879 | origtmp1470;
	assign origtmp59 = in[733] | in[330];
	assign origtmp947 = origtmp950 | origtmp951;
	assign origtmp219 = origtmp218 & origtmp217;
	assign origtmp1545 = in[1310] ^ in[1190];
	assign origtmp2085 = origtmp1310 | origtmp1467;
	assign origtmp293 = origtmp294 ^ origtmp295;
	assign origtmp653 = 1'b1 & origtmp655;
	assign origtmp1482 = in[1391] ^ origtmp1754;
	assign out[78] = origtmp195 | 1'b1;
	assign origtmp252 = ~1'b0;
	assign origtmp123 = in[1034] ^ in[430];
	assign origtmp66 = origtmp68 ^ origtmp68;
	assign out[384] = in[931] & in[318];
	assign origtmp1878 = in[909] & in[918];
	assign origtmp1128 = origtmp1129 ^ origtmp1125;
	assign origtmp761 = origtmp762 ^ in[695];
	assign origtmp899 = 1'b0;
	assign origtmp1443 = origtmp1469 & in[950];
	assign origtmp1195 = origtmp1197 & in[110];
	assign origtmp1608 = in[925] ^ origtmp1403;
	assign origtmp332 = 1'b1 & 1'b1;
	assign origtmp807 = in[169] ^ in[169];
	assign origtmp803 = in[1226] & origtmp805;
	assign out[333] = origtmp833 ^ origtmp831;
	assign out[476] = in[557] ^ in[1239];
	assign origtmp1262 = origtmp1490 | in[1265];
	assign origtmp2073 = origtmp1430 | origtmp1772;
	assign out[395] = origtmp979 ^ in[446];
	assign origtmp1624 = origtmp2117 ^ origtmp1711;
	assign origtmp2217 = origtmp1679 ^ origtmp1824;
	assign origtmp2197 = in[1401] | origtmp2062;
	assign origtmp1791 = origtmp1592 & origtmp1641;
	assign origtmp608 = 1'b0 & origtmp609;
	assign origtmp1152 = 1'b0 ^ 1'b0;
	assign origtmp359 = in[613] ^ 1'b1;
	assign origtmp579 = origtmp578 | in[815];
	assign origtmp73 = origtmp70 & origtmp71;
	assign origtmp1282 = origtmp1817 | origtmp2113;
	assign origtmp2070 = in[62] & in[731];
	assign origtmp977 = origtmp978 | origtmp978;
	assign out[233] = origtmp585 & in[451];
	assign origtmp1368 = origtmp1285 | origtmp1614;
	assign origtmp462 = in[687] | in[715];
	assign origtmp117 = 1'b0;
	assign origtmp1231 = in[610] | in[610];
	assign origtmp1734 = in[1466] ^ in[1065];
	assign origtmp1749 = in[1493] ^ origtmp2130;
	assign out[251] = ~origtmp625;
	assign origtmp2111 = origtmp1603 | origtmp2038;
	assign origtmp836 = ~origtmp835;
	assign origtmp1855 = origtmp1523 & in[712];
	assign out[328] = origtmp816 ^ origtmp814;
	assign origtmp783 = origtmp786 | origtmp784;
	assign out[269] = origtmp669 ^ origtmp672;
	assign origtmp1974 = in[1111] & in[243];
	assign origtmp1954 = origtmp1450 & origtmp2012;
	assign out[487] = origtmp1218 | origtmp1214;
	assign out[102] = origtmp256 & origtmp255;
	assign origtmp154 = origtmp153;
	assign origtmp483 = 1'b0 & origtmp485;
	assign out[173] = origtmp433 | 1'b1;
	assign origtmp1965 = origtmp1522 & origtmp1243;
	assign out[279] = origtmp701 & origtmp703;
	assign origtmp1906 = origtmp1818 & origtmp2222;
	assign origtmp1780 = origtmp1580 ^ in[964];
	assign out[191] = origtmp476 | 1'b0;
	assign out[95] = origtmp240 ^ origtmp241;
	assign origtmp317 = 1'b1 ^ origtmp314;
	assign out[376] = in[478] ^ origtmp929;
	assign out[199] = origtmp500 | origtmp502;
	assign origtmp271 = 1'b1 & origtmp269;
	assign origtmp1346 = origtmp1335 ^ origtmp1673;
	assign origtmp969 = 1'b1 ^ in[704];
	assign origtmp1249 = in[1263] & in[906];
	assign out[162] = in[477] ^ origtmp407;
	assign origtmp370 = in[1387] & in[828];
	assign origtmp1483 = in[324] | in[261];
	assign origtmp28 = in[455] ^ 1'b1;
	assign origtmp1028 = in[1118] & in[1289];
	assign origtmp51 = in[905] ^ in[905];
	assign origtmp694 = in[1021];
	assign origtmp2052 = origtmp1432 ^ origtmp1249;
	assign origtmp2039 = in[865] | in[1058];
	assign out[313] = ~origtmp783;
	assign out[363] = in[468] & in[270];
	assign origtmp1052 = ~1'b0;
	assign origtmp1940 = in[1031] ^ in[1351];
	assign origtmp471 = origtmp473 & origtmp472;
	assign origtmp2100 = origtmp1472 | origtmp1593;
	assign origtmp1747 = origtmp1454 | origtmp1724;
	assign origtmp1220 = origtmp1222 & origtmp1221;
	assign out[491] = in[1141] ^ in[294];
	assign origtmp558 = origtmp557 ^ origtmp559;
	assign origtmp920 = origtmp922 & in[361];
	assign origtmp2022 = origtmp1943 & origtmp1527;
	assign origtmp1913 = origtmp1676 ^ origtmp1375;
	assign origtmp1896 = origtmp1782 ^ origtmp1351;
	assign origtmp1488 = origtmp1349 & origtmp1858;
	assign origtmp1535 = in[409] ^ in[0];
	assign origtmp345 = in[228] ^ 1'b1;
	assign origtmp1138 = ~in[188];
	assign origtmp1442 = origtmp2104 | origtmp2040;
	assign origtmp1342 = origtmp1999 | origtmp1468;
	assign out[309] = in[257] ^ in[399];
	assign origtmp965 = origtmp967 ^ in[1317];
	assign origtmp321 = ~1'b0;
	assign origtmp1980 = in[16] | origtmp1732;
	assign out[71] = origtmp173 | origtmp177;
	assign origtmp1645 = in[820] ^ in[1499];
	assign origtmp482 = 1'b0 ^ origtmp486;
	assign out[237] = origtmp589 & 1'b1;
	assign origtmp580 = origtmp579 | in[815];
	assign origtmp1870 = in[197] | origtmp2138;
	assign origtmp848 = origtmp847 & origtmp846;
	assign out[394] = origtmp977 | 1'b1;
	assign origtmp1347 = in[674] & in[351];
	assign origtmp520 = 1'b1 | in[1172];
	assign origtmp883 = in[286] | in[297];
	assign origtmp1547 = in[835] | origtmp1296;
	assign origtmp2129 = origtmp1401 | origtmp1731;
	assign out[368] = in[386] & in[589];
	assign out[41] = origtmp105 & origtmp105;
	assign origtmp583 = in[775] ^ origtmp581;
	assign origtmp1250 = in[1477] | in[691];
	assign origtmp2013 = origtmp1383 & in[1384];
	assign out[411] = origtmp1009 ^ origtmp1010;
	assign origtmp1703 = origtmp2227 | in[334];
	assign out[132] = in[692] | 1'b1;
	assign origtmp1010 = origtmp1007;
	assign origtmp1851 = in[36] & in[669];
	assign origtmp507 = in[222] & in[922];
	assign origtmp1837 = origtmp1434 ^ in[979];
	assign origtmp240 = 1'b0 | in[1293];
	assign origtmp2135 = in[776] | in[1454];
	assign origtmp835 = 1'b0 & 1'b1;
	assign origtmp1529 = origtmp1761 & origtmp2223;
	assign origtmp1215 = 1'b0 & origtmp1217;
	assign origtmp605 = 1'b1;
	assign origtmp23 = origtmp25 | origtmp26;
	assign origtmp1415 = origtmp1625 | origtmp1791;
	assign origtmp554 = origtmp552 | in[479];
	assign origtmp914 = in[1098];
	assign origtmp2056 = in[80] & in[284];
	assign origtmp181 = in[558] | 1'b0;
	assign out[472] = in[1440] | 1'b1;
	assign origtmp2170 = origtmp1958 | origtmp2160;
	assign origtmp1622 = origtmp1316 & in[30];
	assign origtmp86 = origtmp87 & origtmp90;
	assign out[89] = origtmp222 & 1'b0;
	assign origtmp628 = origtmp630 ^ in[838];
	assign origtmp1478 = in[1273] ^ in[1096];
	assign origtmp1357 = origtmp2194 ^ origtmp1417;
	assign origtmp2156 = origtmp2195 ^ origtmp2198;
	assign origtmp1672 = origtmp1720 & in[313];
	assign origtmp699 = in[757] ^ in[757];
	assign origtmp1307 = origtmp1730 ^ in[864];
	assign origtmp532 = origtmp531 ^ in[203];
	assign origtmp131 = 1'b1 ^ in[953];
	assign origtmp1276 = in[568] & in[1442];
	assign origtmp584 = 1'b1 & origtmp581;
	assign origtmp303 = 1'b1;
	assign out[106] = origtmp267 | in[680];
	assign out[304] = origtmp761 & origtmp761;
	assign origtmp745 = in[235];
	assign origtmp31 = origtmp30 & in[455];
	assign origtmp714 = origtmp715 ^ in[562];
	assign origtmp581 = origtmp582 | 1'b1;
	assign out[441] = origtmp1094 & origtmp1096;
	assign origtmp1424 = origtmp1464 & origtmp1540;
	assign origtmp1605 = in[659] | in[771];
	assign origtmp463 = origtmp465 | 1'b1;
	assign origtmp1521 = origtmp1618 ^ origtmp1405;
	assign origtmp2024 = in[1367] ^ origtmp1485;
	assign origtmp1404 = in[1237] & in[1277];
	assign origtmp850 = ~origtmp852;
	assign out[159] = 1'b1 ^ origtmp397;
	assign origtmp1918 = in[603] & origtmp2237;
	assign origtmp313 = origtmp310 & origtmp309;
	assign origtmp124 = origtmp126;
	assign origtmp189 = 1'b0;
	assign origtmp424 = origtmp423 ^ origtmp422;
	assign origtmp213 = ~1'b0;
	assign origtmp1573 = origtmp1706 | origtmp2165;
	assign origtmp261 = origtmp265 & origtmp265;
	assign origtmp1632 = origtmp1322 ^ origtmp1473;
	assign out[130] = origtmp324 | origtmp324;
	assign out[409] = origtmp1006 ^ origtmp1005;
	assign out[195] = origtmp489 ^ 1'b0;
	assign origtmp348 = origtmp349 ^ origtmp350;
	assign origtmp1673 = in[985] | origtmp1903;
	assign origtmp430 = in[1320] & 1'b0;
	assign origtmp33 = origtmp34 | origtmp32;
	assign origtmp550 = origtmp551 & origtmp549;
	assign out[410] = in[1462] & in[77];
	assign origtmp1419 = origtmp1566 ^ origtmp1571;
	assign origtmp794 = 1'b0;
	assign origtmp384 = in[384];
	assign origtmp1310 = in[429] ^ in[860];
	assign origtmp1146 = origtmp1144 | origtmp1143;
	assign origtmp215 = origtmp216 | origtmp214;
	assign origtmp556 = in[1274] & in[1399];
	assign origtmp856 = in[425] | 1'b1;
	assign out[79] = origtmp196 & 1'b1;
	assign origtmp453 = origtmp452;
	assign out[281] = in[1257] | origtmp708;
	assign origtmp1730 = in[1166] | in[161];
	assign out[31] = in[882];
	assign origtmp2137 = in[145] ^ in[299];
	assign origtmp1746 = origtmp1780 ^ in[1206];
	assign origtmp2248 = in[3] & in[175];
	assign origtmp1126 = in[1216] & 1'b1;
	assign out[415] = origtmp1022 | origtmp1021;
	assign origtmp1530 = origtmp1392 ^ origtmp1877;
	assign origtmp939 = 1'b1 ^ in[551];
	assign origtmp175 = 1'b0 | 1'b1;
	assign origtmp788 = in[310] | 1'b1;
	assign origtmp2062 = origtmp1702 | origtmp1658;
	assign origtmp1013 = origtmp1016 ^ origtmp1014;
	assign origtmp693 = in[1021] & origtmp694;
	assign origtmp2068 = in[861] ^ origtmp1832;
	assign origtmp1205 = origtmp1206 | in[1298];
	assign origtmp141 = in[1051] & in[1051];
	assign origtmp2034 = in[100] | in[1343];
	assign origtmp323 = 1'b0 ^ origtmp321;
	assign origtmp1329 = origtmp1345 & origtmp1948;
	assign origtmp734 = origtmp735 & origtmp731;
	assign origtmp2251 = origtmp2220 ^ origtmp1548;
	assign origtmp814 = origtmp817 ^ in[748];
	assign origtmp1427 = origtmp1827 | in[655];
	assign origtmp1380 = in[484] | origtmp1589;
	assign origtmp470 = origtmp473 & 1'b1;
	assign origtmp108 = 1'b0 ^ origtmp110;
	assign origtmp712 = origtmp710 & origtmp713;
	assign out[316] = origtmp790 | origtmp789;
	assign origtmp1284 = origtmp2084 & in[1192];
	assign origtmp201 = 1'b1 & 1'b0;
	assign origtmp995 = in[47] ^ 1'b0;
	assign origtmp167 = origtmp163 & 1'b0;
	assign origtmp1743 = in[1352] | in[888];
	assign out[298] = in[614] | in[614];
	assign origtmp1201 = ~origtmp1203;
	assign out[348] = origtmp867 & origtmp866;
	assign origtmp510 = 1'b0 | origtmp511;
	assign origtmp1955 = origtmp1493 & origtmp1938;
	assign out[255] = in[503] & origtmp633;
	assign origtmp2253 = in[401] & in[661];
	assign origtmp497 = in[1243] | origtmp495;
	assign origtmp1317 = origtmp1465 ^ origtmp1759;
	assign origtmp1076 = origtmp1075 ^ 1'b0;
	assign origtmp72 = origtmp69 | origtmp73;
	assign origtmp2207 = origtmp1798 | origtmp1539;
	assign origtmp180 = 1'b1 ^ origtmp181;
	assign origtmp1248 = in[1173] ^ origtmp1889;
	assign origtmp1429 = in[211] & in[378];
	assign origtmp797 = 1'b1 & 1'b1;
	assign origtmp2057 = in[955] ^ origtmp1331;
	assign origtmp1280 = in[1283] & in[1375];
	assign origtmp619 = origtmp618 & in[131];
	assign origtmp1397 = in[811] ^ in[21];
	assign origtmp1237 = in[972] | in[474];
	assign out[272] = origtmp679 ^ origtmp680;
	assign origtmp1927 = in[251] & in[460];
	assign origtmp1021 = ~1'b1;
	assign origtmp1150 = 1'b0 | 1'b1;
	assign origtmp417 = in[510] & origtmp415;
	assign origtmp1699 = origtmp1354 & origtmp1549;
	assign origtmp810 = 1'b1 | 1'b0;
	assign origtmp2140 = in[690] | in[215];
	assign out[239] = 1'b1 ^ origtmp597;
	assign origtmp928 = 1'b0 ^ in[354];
	assign out[232] = origtmp583 | origtmp584;
	assign origtmp845 = ~origtmp848;
	assign origtmp1479 = origtmp1555 & in[141];
	assign origtmp1570 = origtmp1833 | origtmp1376;
	assign origtmp1719 = origtmp1687 ^ in[1380];
	assign origtmp50 = origtmp52 ^ in[905];
	assign origtmp1517 = in[1305] ^ origtmp2232;
	assign origtmp1676 = origtmp1635 | origtmp1710;
	assign origtmp765 = origtmp764 | origtmp766;
	assign origtmp1807 = in[424] ^ in[987];
	assign origtmp692 = 1'b0 | 1'b0;
	assign origtmp1843 = origtmp1436 | in[172];
	assign origtmp1630 = origtmp2155 | origtmp1738;
	assign out[152] = in[847] | in[63];
	assign origtmp624 = 1'b0 | origtmp623;
	assign out[311] = 1'b1 | origtmp779;
	assign out[138] = origtmp341 ^ origtmp341;
	assign origtmp948 = 1'b0 ^ origtmp949;
	assign out[332] = origtmp829 ^ origtmp828;
	assign origtmp988 = origtmp989 | origtmp989;
	assign origtmp1299 = origtmp2224 ^ origtmp1851;
	assign origtmp536 = origtmp535 & 1'b1;
	assign origtmp347 = in[1044];
	assign origtmp1585 = origtmp1564 | origtmp1964;
	assign origtmp1773 = in[139] | in[133];
	assign origtmp702 = 1'b1 & in[862];
	assign out[236] = in[1272] & origtmp587;
	assign origtmp654 = origtmp653 & origtmp656;
	assign origtmp1603 = in[1341] ^ in[1406];
	assign out[477] = origtmp1199 ^ in[110];
	assign origtmp2104 = origtmp1488 ^ origtmp1629;
	assign origtmp299 = in[1402] | 1'b1;
	assign origtmp808 = ~origtmp807;
	assign origtmp270 = origtmp268 ^ origtmp271;
	assign origtmp1241 = in[343] | in[711];
	assign out[110] = origtmp278 | 1'b0;
	assign origtmp283 = 1'b1 ^ origtmp281;
	assign origtmp227 = 1'b0;
	assign origtmp1614 = in[8] ^ in[269];
	assign out[0] = origtmp1 | in[626];
	assign origtmp1289 = in[1126] ^ origtmp1516;
	assign out[308] = origtmp773 & origtmp774;
	assign origtmp2035 = origtmp1482 & in[1076];
	assign origtmp1643 = origtmp2187 ^ origtmp1254;
	assign origtmp1803 = origtmp1458 & origtmp1330;
	assign origtmp911 = in[1264] | in[682];
	assign origtmp1664 = origtmp1727 ^ origtmp1448;
	assign out[406] = 1'b1 | origtmp1000;
	assign out[401] = origtmp994 ^ in[1106];
	assign origtmp998 = 1'b0 | origtmp997;
	assign origtmp1111 = ~1'b1;
	assign origtmp546 = 1'b1 | origtmp547;
	assign origtmp1564 = origtmp1763 ^ origtmp1881;
	assign out[153] = origtmp382 | origtmp380;
	assign origtmp894 = in[804] ^ in[1447];
	assign origtmp146 = origtmp143 | in[289];
	assign origtmp1437 = in[254] ^ in[487];
	assign origtmp478 = origtmp481 ^ origtmp481;
	assign origtmp1867 = origtmp2074 | in[359];
	assign origtmp864 = in[148] & in[148];
	assign origtmp1398 = in[143] ^ in[1200];
	assign out[104] = in[851];
	assign origtmp744 = origtmp745 & origtmp743;
	assign origtmp1119 = in[541] & origtmp1115;
	assign origtmp879 = origtmp882 & 1'b0;
	assign origtmp1169 = in[1246] & origtmp1170;
	assign origtmp1826 = origtmp2217 ^ origtmp2170;
	assign origtmp1353 = in[453] | origtmp2216;
	assign origtmp1500 = in[157] | in[974];
	assign origtmp1863 = origtmp1338 | origtmp1935;
	assign origtmp1303 = origtmp1859 | in[11];
	assign origtmp1180 = ~1'b1;
	assign origtmp1168 = in[366] & in[366];
	assign origtmp1463 = origtmp1736 ^ in[402];
	assign origtmp468 = in[501] | in[501];
	assign origtmp2021 = origtmp1916 | origtmp1962;
	assign origtmp1069 = ~origtmp1071;
	assign origtmp963 = 1'b0 & in[230];
	assign origtmp860 = in[138] & 1'b1;
	assign origtmp20 = ~in[87];
	assign out[452] = ~origtmp1130;
	assign origtmp60 = ~origtmp59;
	assign origtmp1300 = in[765] | in[521];
	assign origtmp1122 = origtmp1121 | 1'b0;
	assign origtmp1287 = origtmp1600 & origtmp1767;
	assign origtmp1125 = in[1216] | 1'b0;
	assign origtmp125 = 1'b1 & 1'b1;
	assign origtmp2040 = origtmp2205 & in[729];
	assign out[323] = origtmp802 & origtmp803;
	assign origtmp1852 = origtmp2249 & origtmp1307;
	assign origtmp1019 = ~1'b1;
	assign out[310] = origtmp776 | origtmp778;
	assign origtmp1049 = 1'b1 ^ 1'b1;
	assign origtmp165 = origtmp166 ^ in[320];
	assign origtmp2229 = origtmp1871 | in[1292];
	assign origtmp1629 = origtmp1752 & origtmp2196;
	assign origtmp2001 = origtmp1713 & origtmp2252;
	assign out[124] = origtmp312 | 1'b0;
	assign origtmp781 = in[108] ^ in[502];
	assign origtmp1080 = origtmp1079 | 1'b1;
	assign origtmp1640 = in[774] | in[1496];
	assign origtmp1459 = origtmp1245 ^ in[587];
	assign origtmp1802 = origtmp1582 & in[1382];
	assign origtmp2063 = in[304] & in[586];
	assign origtmp1218 = in[1003] | origtmp1215;
	assign origtmp206 = ~1'b0;
	assign origtmp203 = origtmp201 & origtmp201;
	assign out[3] = origtmp6 ^ origtmp8;
	assign origtmp1050 = 1'b1;
	assign origtmp1788 = in[786] ^ origtmp2179;
	assign out[209] = origtmp517 | in[1218];
	assign origtmp1738 = in[1465] | origtmp1946;
	assign origtmp529 = 1'b0 ^ in[920];
	assign origtmp147 = in[241] ^ origtmp150;
	assign origtmp891 = in[1229] & 1'b0;
	assign origtmp472 = 1'b0 ^ 1'b1;
	assign origtmp1418 = in[1430] & in[1420];
	assign out[96] = 1'b1 ^ origtmp243;
	assign out[372] = origtmp917 | origtmp918;
	assign origtmp1666 = origtmp2246 ^ origtmp1377;
	assign origtmp1510 = in[301] ^ in[193];
	assign origtmp1684 = in[391] & origtmp1524;
	assign origtmp695 = 1'b0 | in[275];
	assign out[458] = origtmp1149 ^ origtmp1148;
	assign origtmp286 = origtmp287 | origtmp284;
	assign origtmp1789 = in[623] ^ in[306];
	assign origtmp2226 = in[588] & in[198];
	assign origtmp1306 = origtmp1491 & origtmp1649;
	assign origtmp780 = 1'b0 & 1'b0;
	assign origtmp429 = in[999] | in[1320];
	assign origtmp407 = in[477] ^ origtmp406;
	assign origtmp221 = in[1062] | in[1437];
	assign out[45] = ~1'b1;
	assign origtmp183 = in[22] ^ 1'b1;
	assign out[183] = 1'b1;
	assign out[26] = 1'b1 ^ origtmp72;
	assign origtmp1403 = origtmp1273 ^ origtmp2058;
	assign origtmp224 = in[1362] & 1'b1;
	assign origtmp427 = in[999] | 1'b1;
	assign origtmp1444 = in[1303] ^ in[296];
	assign out[277] = origtmp698 ^ origtmp696;
	assign origtmp2196 = in[265] | origtmp1489;
	assign origtmp754 = origtmp751;
	assign origtmp1920 = in[673] & in[1043];
	assign origtmp1473 = in[1026] & in[762];
	assign out[252] = origtmp628 | origtmp629;
	assign origtmp1022 = 1'b0;
	assign origtmp1631 = in[1174] & in[620];
	assign out[114] = origtmp288 & 1'b1;
	assign origtmp290 = origtmp291 & 1'b1;
	assign origtmp99 = 1'b1 | 1'b0;
	assign origtmp118 = origtmp115 ^ 1'b1;
	assign origtmp2025 = origtmp1739 | in[741];
	assign origtmp152 = origtmp151;
	assign origtmp1943 = in[345] & in[1093];
	assign origtmp285 = 1'b0;
	assign origtmp1742 = in[1185] | in[1019];
	assign origtmp1236 = ~1'b1;
	assign origtmp812 = in[991] ^ 1'b1;
	assign origtmp1609 = origtmp1945 ^ origtmp1995;
	assign out[457] = 1'b1 & origtmp1147;
	assign out[221] = origtmp553 & origtmp555;
	assign origtmp1519 = in[1235] & in[1389];
	assign origtmp2216 = origtmp1586 & in[262];
	assign origtmp1895 = origtmp1758 & origtmp2218;
	assign origtmp433 = origtmp435;
	assign out[156] = origtmp389 & origtmp386;
	assign origtmp1889 = in[758] ^ in[752];
	assign out[342] = origtmp853 ^ origtmp855;
	assign out[74] = origtmp184 & in[22];
	assign out[350] = origtmp871 ^ origtmp871;
	assign origtmp853 = origtmp854 ^ origtmp854;
	assign origtmp2122 = in[58] ^ origtmp2197;
	assign origtmp1994 = origtmp1662 ^ origtmp2128;
	assign origtmp35 = 1'b0;
	assign origtmp2106 = in[998] & origtmp1503;
	assign origtmp1827 = origtmp1801 & origtmp1869;
	assign out[349] = origtmp868 ^ origtmp869;
	assign origtmp1933 = origtmp1399 ^ in[967];
	assign origtmp844 = 1'b1 | 1'b1;
	assign origtmp668 = in[632] | in[495];
	assign origtmp1183 = origtmp1187 & 1'b1;
	assign origtmp1043 = origtmp1042;
	assign out[77] = in[439] & origtmp190;
	assign origtmp1273 = in[713] ^ in[49];
	assign out[68] = ~1'b1;
	assign origtmp2209 = origtmp1803 | in[379];
	assign origtmp2041 = in[1102] | in[271];
	assign origtmp102 = origtmp103 | origtmp100;
	assign origtmp527 = ~origtmp526;
	assign origtmp2220 = origtmp1483 & origtmp1795;
	assign out[178] = 1'b0;
	assign origtmp431 = origtmp429 ^ origtmp430;
	assign origtmp1064 = in[726] ^ in[938];
	assign origtmp728 = 1'b1 ^ in[388];
	assign origtmp75 = origtmp74 ^ origtmp74;
	assign origtmp295 = 1'b1;
	assign origtmp627 = 1'b0 ^ 1'b1;
	assign origtmp1266 = origtmp1334 & origtmp1919;
	assign origtmp972 = in[567] | origtmp971;
	assign origtmp392 = ~origtmp391;
	assign origtmp1593 = in[635] | origtmp2174;
	assign origtmp1359 = in[993] & in[658];
	assign origtmp1063 = 1'b1 | in[369];
	assign out[179] = origtmp445 ^ origtmp443;
	assign origtmp631 = in[1479] & in[1479];
	assign origtmp1323 = in[877] ^ in[990];
	assign origtmp222 = in[647] | in[574];
	assign origtmp1833 = origtmp1927 & origtmp1921;
	assign origtmp2240 = in[50] & in[517];
	assign origtmp2238 = origtmp1846 & in[1251];
	assign origtmp375 = 1'b0 & in[1002];
	assign origtmp404 = 1'b1;
	assign origtmp1198 = in[110] ^ in[660];
	assign out[157] = origtmp394 ^ origtmp395;
	assign out[91] = origtmp227;
	assign origtmp726 = in[388] | 1'b1;
	assign origtmp1989 = origtmp2158 ^ origtmp2006;
	assign origtmp1014 = origtmp1012 & origtmp1012;
	assign origtmp1656 = in[292] | origtmp1427;
	assign origtmp1924 = in[639] & origtmp2193;
	assign out[339] = origtmp844 | origtmp845;
	assign origtmp1200 = ~1'b1;
	assign origtmp226 = origtmp223 & in[1362];
	assign origtmp1430 = in[736] ^ in[170];
	assign origtmp1618 = in[844] ^ origtmp1444;
	assign out[247] = origtmp616 & origtmp614;
	assign origtmp1950 = in[1045] | in[370];
	assign origtmp1085 = 1'b0;
	assign origtmp1277 = in[797] & in[932];
	assign origtmp1612 = in[686] | in[104];
	assign origtmp1650 = origtmp1563 ^ in[935];
	assign origtmp533 = in[1415] & origtmp534;
	assign origtmp199 = in[350] & 1'b0;
	assign origtmp809 = 1'b1 & 1'b0;
	assign origtmp612 = in[258] ^ in[650];
	assign origtmp1321 = in[1079] & in[556];
	assign origtmp2136 = origtmp2002 | origtmp1888;
	assign out[48] = origtmp118 | origtmp116;
	assign origtmp659 = 1'b0 ^ origtmp658;
	assign origtmp1056 = 1'b0 | origtmp1052;
	assign origtmp1039 = in[122] | 1'b0;
	assign out[118] = 1'b1 | origtmp293;
	assign origtmp1982 = in[1146] ^ origtmp2009;
	assign origtmp2003 = in[410] ^ in[789];
	assign origtmp818 = origtmp815 & 1'b0;
	assign origtmp1537 = in[309] & origtmp1714;
	assign out[217] = origtmp538 | 1'b0;
	assign origtmp1234 = in[136] & 1'b1;
	assign origtmp231 = ~1'b0;
	assign origtmp1579 = in[1432] | origtmp1255;
	assign origtmp316 = in[98] & origtmp315;
	assign origtmp1764 = in[1001] & origtmp1944;
	assign origtmp179 = 1'b1 ^ origtmp180;
	assign origtmp2223 = in[1448] & in[1459];
	assign origtmp93 = in[796];
	assign origtmp1588 = in[73] & in[1327];
	assign out[116] = in[1061] ^ in[1168];
	assign origtmp1147 = in[1480] ^ in[1480];
	assign origtmp381 = in[1315] ^ 1'b0;
	assign origtmp1191 = origtmp1190;
	assign origtmp1105 = 1'b0;
	assign origtmp1963 = in[1356] | origtmp1863;
	assign origtmp15 = origtmp13 & origtmp12;
	assign origtmp719 = 1'b1;
	assign origtmp1005 = origtmp1004 & 1'b1;
	assign origtmp136 = ~in[1032];
	assign origtmp78 = origtmp80 | origtmp79;
	assign origtmp2233 = origtmp1917 & in[1135];
	assign out[244] = 1'b0;
	assign origtmp2038 = in[1040] | in[699];
	assign origtmp986 = origtmp985 ^ origtmp985;
	assign origtmp2096 = origtmp1451 ^ in[1470];
	assign origtmp589 = origtmp588 ^ origtmp588;
	assign origtmp143 = origtmp142 & in[289];
	assign origtmp1061 = 1'b0;
	assign out[225] = origtmp567;
	assign origtmp820 = 1'b0 | in[210];
	assign origtmp679 = origtmp678 & 1'b1;
	assign out[20] = in[1101] | origtmp53;
	assign origtmp406 = 1'b0 ^ origtmp405;
	assign origtmp1256 = in[1476] & in[238];
	assign origtmp542 = origtmp545 | origtmp541;
	assign origtmp1669 = origtmp1876 & origtmp1590;
	assign origtmp645 = 1'b0;
	assign origtmp1623 = in[389] & in[1256];
	assign origtmp1596 = in[209] | in[1122];
	assign origtmp1725 = in[525] & in[23];
	assign origtmp437 = origtmp438 | 1'b0;
	assign origtmp19 = origtmp18 & origtmp18;
	assign origtmp1713 = origtmp1342 & origtmp1312;
	assign origtmp1090 = 1'b0 | origtmp1087;
	assign origtmp1041 = origtmp1039 & origtmp1040;
	assign origtmp1245 = origtmp1744 ^ in[744];
	assign origtmp385 = origtmp384 ^ 1'b0;
	assign origtmp731 = origtmp733;
	assign origtmp936 = 1'b0 & in[1498];
	assign origtmp207 = origtmp206;
	assign origtmp2202 = origtmp2000 ^ in[126];
	assign origtmp502 = origtmp501;
	assign out[360] = ~1'b0;
	assign origtmp1864 = origtmp2253 ^ in[832];
	assign origtmp1836 = in[937] ^ in[592];
	assign origtmp2249 = origtmp1550 & origtmp1616;
	assign origtmp717 = 1'b0 | 1'b0;
	assign origtmp1655 = origtmp1960 & in[353];
	assign origtmp1987 = origtmp1779 | in[770];
	assign origtmp2049 = in[109] ^ in[805];
	assign origtmp576 = ~1'b1;
	assign origtmp1528 = in[40] & in[154];
	assign origtmp1335 = origtmp2069 & in[1266];
	assign origtmp354 = 1'b1 ^ 1'b1;
	assign origtmp681 = 1'b1 ^ 1'b0;
	assign origtmp528 = ~in[1414];
	assign origtmp1409 = origtmp1284 ^ origtmp1703;
	assign origtmp925 = in[478] | in[478];
	assign origtmp964 = in[105] | 1'b0;
	assign origtmp2230 = origtmp1637 & origtmp1353;
	assign origtmp1541 = in[969] ^ origtmp2065;
	assign origtmp1838 = origtmp2036 & origtmp1274;
	assign origtmp191 = origtmp194 & origtmp194;
	assign origtmp521 = 1'b0 & in[444];
	assign origtmp300 = origtmp301 & origtmp299;
	assign origtmp824 = 1'b0 ^ 1'b0;
	assign origtmp971 = in[704] & in[567];
	assign out[35] = origtmp95 | origtmp95;
	assign origtmp1748 = origtmp1587 & in[373];
	assign origtmp30 = origtmp28 | 1'b1;
	assign origtmp825 = origtmp827 | in[1458];
	assign origtmp1999 = in[1259] | in[514];
	assign origtmp614 = origtmp613 & in[650];
	assign origtmp1309 = in[372] ^ origtmp2207;
	assign origtmp1681 = origtmp2124 ^ in[666];
	assign origtmp1449 = in[1] & in[1485];
	assign origtmp867 = in[1429] | in[148];
	assign origtmp1894 = origtmp2017 & origtmp1769;
	assign out[388] = origtmp958 ^ origtmp957;
	assign origtmp1475 = in[1212] ^ in[897];
	assign origtmp1468 = origtmp2011 | origtmp1907;
	assign origtmp2192 = origtmp2061 & origtmp1913;
	assign origtmp328 = 1'b0 ^ 1'b0;
	assign origtmp200 = 1'b0 | 1'b0;
	assign origtmp2204 = origtmp2086 & origtmp1678;
	assign origtmp195 = origtmp191 ^ origtmp193;
	assign origtmp2000 = origtmp1682 ^ in[293];
	assign origtmp1910 = in[911] & in[196];
	assign out[317] = in[481] | origtmp792;
	assign origtmp1062 = in[1423] & in[369];
	assign origtmp846 = 1'b0;
	assign origtmp1811 = in[327] ^ in[158];
	assign origtmp357 = in[390] ^ origtmp354;
	assign out[291] = origtmp739 ^ origtmp736;
	assign origtmp505 = 1'b1 | in[822];
	assign origtmp700 = in[757] | in[757];
	assign origtmp2006 = origtmp1605 ^ origtmp2202;
	assign out[396] = 1'b0 & origtmp980;
	assign out[321] = in[853] & origtmp796;
	assign out[354] = origtmp884;
	assign out[61] = in[812] ^ origtmp152;
	assign origtmp898 = 1'b0 & 1'b1;
	assign out[108] = origtmp277 & origtmp273;
	assign origtmp672 = origtmp671 & origtmp670;
	assign origtmp2134 = in[1070] ^ in[1066];
	assign origtmp1816 = origtmp2256 & origtmp2136;
	assign origtmp560 = 1'b1 ^ in[942];
	assign origtmp1214 = origtmp1216 | 1'b1;
	assign origtmp577 = 1'b1;
	assign origtmp1226 = 1'b1 | 1'b1;
	assign origtmp194 = origtmp192 ^ 1'b1;
	assign out[230] = origtmp577 ^ origtmp577;
	assign out[497] = origtmp1235 & origtmp1236;
	assign out[456] = origtmp1146 | in[328];
	assign origtmp1985 = in[1326] ^ in[1017];
	assign origtmp140 = ~in[1018];
	assign origtmp1354 = in[187] | origtmp1853;
	assign origtmp1182 = ~1'b0;
	assign out[365] = in[829] ^ in[1138];
	assign origtmp1544 = origtmp1972 & in[594];
	assign origtmp1003 = 1'b0 ^ 1'b1;
	assign origtmp1078 = ~1'b0;
	assign origtmp1657 = origtmp1987 | in[530];
	assign origtmp1453 = in[509] & in[978];
	assign origtmp119 = origtmp120 ^ origtmp122;
	assign origtmp1425 = origtmp2200 & origtmp2228;
	assign origtmp1759 = origtmp1965 & origtmp1433;
	assign origtmp21 = origtmp17 ^ in[87];
	assign origtmp541 = origtmp543 | origtmp543;
	assign out[444] = origtmp1103 ^ in[1047];
	assign origtmp1455 = origtmp1404 & in[1438];
	assign out[429] = origtmp1065 & origtmp1067;
	assign origtmp122 = 1'b0 & in[83];
	assign origtmp1969 = in[1008] ^ in[12];
	assign origtmp632 = 1'b0;
	assign origtmp177 = origtmp175 ^ origtmp174;
	assign origtmp1938 = in[1262] | in[416];
	assign origtmp908 = origtmp907 ^ in[316];
	assign out[421] = in[1311] | origtmp1041;
	assign origtmp372 = origtmp374 | origtmp374;
	assign origtmp150 = origtmp149;
	assign origtmp421 = ~1'b1;
	assign origtmp667 = 1'b0 & 1'b0;
	assign origtmp616 = 1'b1 ^ 1'b1;
	assign origtmp1098 = origtmp1099 | in[636];
	assign out[470] = origtmp1178 ^ origtmp1182;
	assign origtmp343 = in[228] ^ origtmp344;
	assign origtmp109 = 1'b1 | origtmp110;
	assign origtmp1520 = in[570] & in[195];
	assign origtmp1318 = in[997] | in[1377];
	assign out[392] = origtmp969 & origtmp970;
	assign out[399] = origtmp990 | 1'b0;
	assign origtmp1474 = in[664] | in[102];
	assign origtmp1704 = origtmp2054 & in[867];
	assign origtmp353 = 1'b0 & origtmp351;
	assign origtmp2160 = origtmp1326 ^ origtmp1978;
	assign origtmp1456 = in[1209] ^ origtmp1988;
	assign out[471] = 1'b1 | origtmp1186;
	assign origtmp690 = 1'b0;
	assign origtmp428 = origtmp427 ^ origtmp429;
	assign origtmp2108 = origtmp1882 | origtmp2078;
	assign out[329] = origtmp822 & origtmp823;
	assign origtmp2212 = origtmp1844 ^ origtmp2177;
	assign origtmp2210 = in[1488] | origtmp2153;
	assign origtmp352 = 1'b0 ^ origtmp351;
	assign origtmp488 = origtmp487 ^ origtmp490;
	assign origtmp1893 = origtmp2067 & origtmp1396;
	assign origtmp2144 = in[628] ^ origtmp1839;
	assign origtmp1663 = origtmp1511 | origtmp2001;
	assign origtmp2060 = origtmp1866 | origtmp1954;
	assign origtmp1683 = in[1351] ^ origtmp1947;
	assign out[271] = 1'b0 ^ origtmp677;
	assign origtmp1620 = origtmp1387 | origtmp1319;
	assign out[227] = in[1060] & in[411];
	assign origtmp1511 = origtmp1313 & origtmp1819;
	assign out[382] = origtmp941 & 1'b1;
	assign origtmp1744 = in[1308] | in[565];
	assign origtmp650 = 1'b1 ^ origtmp652;
endmodule

module tb();
    reg[499:0] results[1];
    reg[1499:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%1500b]", data[0]);
        #1
        $display("results = [%500b]", results[0]);
        $writememb("results.txt", results);
    end
endmodule

