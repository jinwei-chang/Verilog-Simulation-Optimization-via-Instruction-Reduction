module dut (out, in);
	output[9:0] out;
	input[29:0] in;
	wire origtmp1;
	wire origtmp2;
	wire origtmp3;
	wire origtmp4;
	wire origtmp5;
	wire origtmp6;
	wire origtmp7;
	wire origtmp8;
	wire origtmp9;
	wire origtmp10;
	wire origtmp11;
	wire origtmp12;
	wire origtmp13;
	wire origtmp14;
	wire origtmp15;
	wire origtmp16;
	wire origtmp17;
	wire origtmp18;
	wire origtmp19;
	wire origtmp20;
	wire origtmp21;
	wire origtmp22;
	wire origtmp23;
	wire origtmp24;
	wire origtmp25;
	wire origtmp26;
	wire origtmp27;
	wire origtmp28;
	wire origtmp29;
	wire origtmp30;
	wire origtmp31;
	wire origtmp32;
	wire origtmp33;
	wire origtmp34;
	wire origtmp35;
	wire origtmp36;
	assign out[0] = origtmp1 | origtmp24;
	assign origtmp1 = origtmp2 | origtmp21;
	assign origtmp2 = origtmp3 | origtmp18;
	assign origtmp3 = origtmp4 | origtmp15;
	assign origtmp4 = origtmp5 | origtmp9;
	assign origtmp5 = in[17] & origtmp6;
	assign origtmp6 = origtmp7 | in[25];
	assign origtmp7 = in[9] & origtmp8;
	assign origtmp8 = in[6] & in[27];
	assign origtmp9 = origtmp10 ^ origtmp14;
	assign origtmp10 = origtmp11 | origtmp12;
	assign origtmp11 = in[7] | in[26];
	assign origtmp12 = origtmp13 & in[10];
	assign origtmp13 = in[5] & in[13];
	assign origtmp14 = in[8] | in[2];
	assign origtmp15 = in[19] ^ origtmp16;
	assign origtmp16 = origtmp17 & in[4];
	assign origtmp17 = in[21] ^ in[12];
	assign origtmp18 = origtmp19 & origtmp20;
	assign origtmp19 = in[24] & in[23];
	assign origtmp20 = in[14] | in[20];
	assign origtmp21 = origtmp22 & origtmp23;
	assign origtmp22 = in[3] | in[1];
	assign origtmp23 = in[15] ^ in[16];
	assign origtmp24 = 1'b1 | origtmp25;
	assign origtmp25 = origtmp26 | origtmp30;
	assign origtmp26 = origtmp27 & origtmp28;
	assign origtmp27 = in[11] | in[24];
	assign origtmp28 = in[22] & origtmp29;
	assign origtmp29 = in[0] | in[18];
	assign origtmp30 = in[24] | origtmp31;
	assign origtmp31 = in[24] & in[21];
	assign out[1] = origtmp32 ^ in[28];
	assign origtmp32 = 1'b1 & 1'b0;
	assign out[2] = 1'b1 & 1'b0;
	assign out[3] = origtmp33;
	assign origtmp33 = 1'b1 & 1'b0;
	assign out[4] = 1'b0 ^ 1'b0;
	assign out[5] = 1'b1;
	assign out[6] = 1'b1 | origtmp34;
	assign origtmp34 = ~1'b0;
	assign out[7] = 1'b0 | origtmp35;
	assign origtmp35 = 1'b0;
	assign out[8] = 1'b0;
	assign out[9] = 1'b1 & origtmp36;
	assign origtmp36 = in[29] | 1'b0;
endmodule

module tb();
    reg[9:0] results[1];
    reg[29:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%30b]", data[0]);
        #1
        $display("results = [%10b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
