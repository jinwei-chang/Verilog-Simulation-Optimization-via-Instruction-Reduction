module dut (out, in);
	output[6:0] out;
	input[35:0] in;
	wire xformtmp15;
	assign xformtmp15 = ~in[27];
	wire xformtmp38;
	assign xformtmp38 = in[29] & xformtmp15;
	wire xformtmp37;
	assign xformtmp37 = ~xformtmp38;
	wire xformtmp17;
	assign xformtmp17 = ~in[31];
	wire xformtmp40;
	assign xformtmp40 = in[33] & xformtmp17;
	wire xformtmp39;
	assign xformtmp39 = ~xformtmp40;
	wire xformtmp74;
	assign xformtmp74 = xformtmp37 & xformtmp39;
	wire xformtmp13;
	assign xformtmp13 = ~in[23];
	wire xformtmp36;
	assign xformtmp36 = in[25] & xformtmp13;
	wire xformtmp35;
	assign xformtmp35 = ~xformtmp36;
	wire xformtmp75;
	assign xformtmp75 = xformtmp74 & xformtmp35;
	wire xformtmp11;
	assign xformtmp11 = ~in[19];
	wire xformtmp34;
	assign xformtmp34 = in[21] & xformtmp11;
	wire xformtmp33;
	assign xformtmp33 = ~xformtmp34;
	wire xformtmp76;
	assign xformtmp76 = xformtmp75 & xformtmp33;
	wire xformtmp9;
	assign xformtmp9 = ~in[15];
	wire xformtmp32;
	assign xformtmp32 = in[17] & xformtmp9;
	wire xformtmp31;
	assign xformtmp31 = ~xformtmp32;
	wire xformtmp77;
	assign xformtmp77 = xformtmp76 & xformtmp31;
	wire xformtmp7;
	assign xformtmp7 = ~in[11];
	wire xformtmp30;
	assign xformtmp30 = in[13] & xformtmp7;
	wire xformtmp29;
	assign xformtmp29 = ~xformtmp30;
	wire xformtmp78;
	assign xformtmp78 = xformtmp77 & xformtmp29;
	wire xformtmp5;
	assign xformtmp5 = ~in[7];
	wire xformtmp28;
	assign xformtmp28 = in[9] & xformtmp5;
	wire xformtmp27;
	assign xformtmp27 = ~xformtmp28;
	wire xformtmp79;
	assign xformtmp79 = xformtmp78 & xformtmp27;
	wire xformtmp3;
	assign xformtmp3 = ~in[3];
	wire xformtmp26;
	assign xformtmp26 = in[5] & xformtmp3;
	wire xformtmp25;
	assign xformtmp25 = ~xformtmp26;
	wire xformtmp80;
	assign xformtmp80 = xformtmp79 & xformtmp25;
	wire xformtmp1;
	assign xformtmp1 = ~in[0];
	wire xformtmp20;
	assign xformtmp20 = in[1] & xformtmp1;
	wire xformtmp19;
	assign xformtmp19 = ~xformtmp20;
	wire xformtmp73;
	assign xformtmp73 = xformtmp80 & xformtmp19;
	assign out[0] = ~xformtmp73;
	wire xformtmp81;
	assign xformtmp81 = ~xformtmp73;
	wire xformtmp94;
	assign xformtmp94 = xformtmp81 ^ xformtmp37;
	wire xformtmp16;
	assign xformtmp16 = ~in[29];
	wire xformtmp66;
	assign xformtmp66 = in[30] | xformtmp16;
	wire xformtmp65;
	assign xformtmp65 = ~xformtmp66;
	wire xformtmp127;
	assign xformtmp127 = xformtmp94 & xformtmp65;
	wire xformtmp126;
	assign xformtmp126 = ~xformtmp127;
	wire xformtmp97;
	assign xformtmp97 = xformtmp81 ^ xformtmp39;
	wire xformtmp18;
	assign xformtmp18 = ~in[33];
	wire xformtmp70;
	assign xformtmp70 = in[34] | xformtmp18;
	wire xformtmp69;
	assign xformtmp69 = ~xformtmp70;
	wire xformtmp129;
	assign xformtmp129 = xformtmp97 & xformtmp69;
	wire xformtmp128;
	assign xformtmp128 = ~xformtmp129;
	wire xformtmp147;
	assign xformtmp147 = xformtmp126 & xformtmp128;
	wire xformtmp91;
	assign xformtmp91 = xformtmp81 ^ xformtmp35;
	wire xformtmp14;
	assign xformtmp14 = ~in[25];
	wire xformtmp62;
	assign xformtmp62 = in[26] | xformtmp14;
	wire xformtmp61;
	assign xformtmp61 = ~xformtmp62;
	wire xformtmp125;
	assign xformtmp125 = xformtmp91 & xformtmp61;
	wire xformtmp124;
	assign xformtmp124 = ~xformtmp125;
	wire xformtmp148;
	assign xformtmp148 = xformtmp147 & xformtmp124;
	wire xformtmp88;
	assign xformtmp88 = xformtmp81 ^ xformtmp33;
	wire xformtmp12;
	assign xformtmp12 = ~in[21];
	wire xformtmp58;
	assign xformtmp58 = in[22] | xformtmp12;
	wire xformtmp57;
	assign xformtmp57 = ~xformtmp58;
	wire xformtmp123;
	assign xformtmp123 = xformtmp88 & xformtmp57;
	wire xformtmp122;
	assign xformtmp122 = ~xformtmp123;
	wire xformtmp149;
	assign xformtmp149 = xformtmp148 & xformtmp122;
	wire xformtmp87;
	assign xformtmp87 = xformtmp81 ^ xformtmp31;
	wire xformtmp10;
	assign xformtmp10 = ~in[17];
	wire xformtmp54;
	assign xformtmp54 = in[18] | xformtmp10;
	wire xformtmp53;
	assign xformtmp53 = ~xformtmp54;
	wire xformtmp121;
	assign xformtmp121 = xformtmp87 & xformtmp53;
	wire xformtmp120;
	assign xformtmp120 = ~xformtmp121;
	wire xformtmp150;
	assign xformtmp150 = xformtmp149 & xformtmp120;
	wire xformtmp86;
	assign xformtmp86 = xformtmp81 ^ xformtmp29;
	wire xformtmp8;
	assign xformtmp8 = ~in[13];
	wire xformtmp50;
	assign xformtmp50 = in[14] | xformtmp8;
	wire xformtmp49;
	assign xformtmp49 = ~xformtmp50;
	wire xformtmp119;
	assign xformtmp119 = xformtmp86 & xformtmp49;
	wire xformtmp118;
	assign xformtmp118 = ~xformtmp119;
	wire xformtmp151;
	assign xformtmp151 = xformtmp150 & xformtmp118;
	wire xformtmp85;
	assign xformtmp85 = xformtmp81 ^ xformtmp27;
	wire xformtmp6;
	assign xformtmp6 = ~in[9];
	wire xformtmp46;
	assign xformtmp46 = in[10] | xformtmp6;
	wire xformtmp45;
	assign xformtmp45 = ~xformtmp46;
	wire xformtmp117;
	assign xformtmp117 = xformtmp85 & xformtmp45;
	wire xformtmp116;
	assign xformtmp116 = ~xformtmp117;
	wire xformtmp152;
	assign xformtmp152 = xformtmp151 & xformtmp116;
	wire xformtmp84;
	assign xformtmp84 = xformtmp81 ^ xformtmp25;
	wire xformtmp4;
	assign xformtmp4 = ~in[5];
	wire xformtmp42;
	assign xformtmp42 = in[6] | xformtmp4;
	wire xformtmp41;
	assign xformtmp41 = ~xformtmp42;
	wire xformtmp115;
	assign xformtmp115 = xformtmp84 & xformtmp41;
	wire xformtmp114;
	assign xformtmp114 = ~xformtmp115;
	wire xformtmp153;
	assign xformtmp153 = xformtmp152 & xformtmp114;
	wire xformtmp83;
	assign xformtmp83 = xformtmp81 ^ xformtmp19;
	wire xformtmp2;
	assign xformtmp2 = ~in[1];
	wire xformtmp22;
	assign xformtmp22 = in[2] | xformtmp2;
	wire xformtmp21;
	assign xformtmp21 = ~xformtmp22;
	wire xformtmp111;
	assign xformtmp111 = xformtmp83 & xformtmp21;
	wire xformtmp110;
	assign xformtmp110 = ~xformtmp111;
	wire xformtmp146;
	assign xformtmp146 = xformtmp153 & xformtmp110;
	assign out[1] = ~xformtmp146;
	wire xformtmp163;
	assign xformtmp163 = ~xformtmp146;
	wire xformtmp180;
	assign xformtmp180 = xformtmp163 ^ xformtmp126;
	wire xformtmp68;
	assign xformtmp68 = in[32] | xformtmp16;
	wire xformtmp67;
	assign xformtmp67 = ~xformtmp68;
	wire xformtmp143;
	assign xformtmp143 = xformtmp94 & xformtmp67;
	wire xformtmp207;
	assign xformtmp207 = xformtmp180 & xformtmp143;
	wire xformtmp206;
	assign xformtmp206 = ~xformtmp207;
	wire xformtmp183;
	assign xformtmp183 = xformtmp163 ^ xformtmp128;
	wire xformtmp72;
	assign xformtmp72 = in[35] | xformtmp18;
	wire xformtmp71;
	assign xformtmp71 = ~xformtmp72;
	wire xformtmp145;
	assign xformtmp145 = xformtmp97 & xformtmp71;
	wire xformtmp209;
	assign xformtmp209 = xformtmp183 & xformtmp145;
	wire xformtmp208;
	assign xformtmp208 = ~xformtmp209;
	wire xformtmp211;
	assign xformtmp211 = xformtmp206 & xformtmp208;
	wire xformtmp177;
	assign xformtmp177 = xformtmp163 ^ xformtmp124;
	wire xformtmp64;
	assign xformtmp64 = in[28] | xformtmp14;
	wire xformtmp63;
	assign xformtmp63 = ~xformtmp64;
	wire xformtmp141;
	assign xformtmp141 = xformtmp91 & xformtmp63;
	wire xformtmp205;
	assign xformtmp205 = xformtmp177 & xformtmp141;
	wire xformtmp204;
	assign xformtmp204 = ~xformtmp205;
	wire xformtmp212;
	assign xformtmp212 = xformtmp211 & xformtmp204;
	wire xformtmp174;
	assign xformtmp174 = xformtmp163 ^ xformtmp122;
	wire xformtmp60;
	assign xformtmp60 = in[24] | xformtmp12;
	wire xformtmp59;
	assign xformtmp59 = ~xformtmp60;
	wire xformtmp139;
	assign xformtmp139 = xformtmp88 & xformtmp59;
	wire xformtmp203;
	assign xformtmp203 = xformtmp174 & xformtmp139;
	wire xformtmp202;
	assign xformtmp202 = ~xformtmp203;
	wire xformtmp213;
	assign xformtmp213 = xformtmp212 & xformtmp202;
	wire xformtmp171;
	assign xformtmp171 = xformtmp163 ^ xformtmp120;
	wire xformtmp56;
	assign xformtmp56 = in[20] | xformtmp10;
	wire xformtmp55;
	assign xformtmp55 = ~xformtmp56;
	wire xformtmp137;
	assign xformtmp137 = xformtmp87 & xformtmp55;
	wire xformtmp201;
	assign xformtmp201 = xformtmp171 & xformtmp137;
	wire xformtmp200;
	assign xformtmp200 = ~xformtmp201;
	wire xformtmp214;
	assign xformtmp214 = xformtmp213 & xformtmp200;
	wire xformtmp168;
	assign xformtmp168 = xformtmp163 ^ xformtmp118;
	wire xformtmp52;
	assign xformtmp52 = in[16] | xformtmp8;
	wire xformtmp51;
	assign xformtmp51 = ~xformtmp52;
	wire xformtmp135;
	assign xformtmp135 = xformtmp86 & xformtmp51;
	wire xformtmp199;
	assign xformtmp199 = xformtmp168 & xformtmp135;
	wire xformtmp198;
	assign xformtmp198 = ~xformtmp199;
	wire xformtmp215;
	assign xformtmp215 = xformtmp214 & xformtmp198;
	wire xformtmp167;
	assign xformtmp167 = xformtmp163 ^ xformtmp116;
	wire xformtmp48;
	assign xformtmp48 = in[12] | xformtmp6;
	wire xformtmp47;
	assign xformtmp47 = ~xformtmp48;
	wire xformtmp133;
	assign xformtmp133 = xformtmp85 & xformtmp47;
	wire xformtmp197;
	assign xformtmp197 = xformtmp167 & xformtmp133;
	wire xformtmp196;
	assign xformtmp196 = ~xformtmp197;
	wire xformtmp216;
	assign xformtmp216 = xformtmp215 & xformtmp196;
	wire xformtmp166;
	assign xformtmp166 = xformtmp163 ^ xformtmp114;
	wire xformtmp44;
	assign xformtmp44 = in[8] | xformtmp4;
	wire xformtmp43;
	assign xformtmp43 = ~xformtmp44;
	wire xformtmp131;
	assign xformtmp131 = xformtmp84 & xformtmp43;
	wire xformtmp195;
	assign xformtmp195 = xformtmp166 & xformtmp131;
	wire xformtmp194;
	assign xformtmp194 = ~xformtmp195;
	wire xformtmp217;
	assign xformtmp217 = xformtmp216 & xformtmp194;
	wire xformtmp165;
	assign xformtmp165 = xformtmp163 ^ xformtmp110;
	wire xformtmp24;
	assign xformtmp24 = in[4] | xformtmp2;
	wire xformtmp23;
	assign xformtmp23 = ~xformtmp24;
	wire xformtmp113;
	assign xformtmp113 = xformtmp83 & xformtmp23;
	wire xformtmp193;
	assign xformtmp193 = xformtmp165 & xformtmp113;
	wire xformtmp192;
	assign xformtmp192 = ~xformtmp193;
	wire xformtmp210;
	assign xformtmp210 = xformtmp217 & xformtmp192;
	assign out[2] = ~xformtmp210;
	wire xformtmp164;
	assign xformtmp164 = ~xformtmp146;
	wire xformtmp170;
	assign xformtmp170 = in[2] & xformtmp164;
	wire xformtmp169;
	assign xformtmp169 = ~xformtmp170;
	wire xformtmp218;
	assign xformtmp218 = ~xformtmp210;
	wire xformtmp220;
	assign xformtmp220 = in[4] & xformtmp218;
	wire xformtmp219;
	assign xformtmp219 = ~xformtmp220;
	wire xformtmp238;
	assign xformtmp238 = xformtmp169 & xformtmp219;
	wire xformtmp82;
	assign xformtmp82 = ~xformtmp73;
	wire xformtmp90;
	assign xformtmp90 = in[0] & xformtmp82;
	wire xformtmp89;
	assign xformtmp89 = ~xformtmp90;
	wire xformtmp239;
	assign xformtmp239 = xformtmp238 & xformtmp89;
	wire xformtmp240;
	assign xformtmp240 = in[1] & xformtmp239;
	wire xformtmp234;
	assign xformtmp234 = in[32] & xformtmp218;
	wire xformtmp233;
	assign xformtmp233 = ~xformtmp234;
	wire xformtmp266;
	assign xformtmp266 = in[29] & xformtmp233;
	wire xformtmp189;
	assign xformtmp189 = in[30] & xformtmp164;
	wire xformtmp188;
	assign xformtmp188 = ~xformtmp189;
	wire xformtmp267;
	assign xformtmp267 = xformtmp266 & xformtmp188;
	wire xformtmp107;
	assign xformtmp107 = in[27] & xformtmp82;
	wire xformtmp106;
	assign xformtmp106 = ~xformtmp107;
	wire xformtmp268;
	assign xformtmp268 = xformtmp267 & xformtmp106;
	wire xformtmp265;
	assign xformtmp265 = ~xformtmp268;
	wire xformtmp236;
	assign xformtmp236 = in[35] & xformtmp218;
	wire xformtmp235;
	assign xformtmp235 = ~xformtmp236;
	wire xformtmp270;
	assign xformtmp270 = in[33] & xformtmp235;
	wire xformtmp191;
	assign xformtmp191 = in[34] & xformtmp164;
	wire xformtmp190;
	assign xformtmp190 = ~xformtmp191;
	wire xformtmp271;
	assign xformtmp271 = xformtmp270 & xformtmp190;
	wire xformtmp109;
	assign xformtmp109 = in[31] & xformtmp82;
	wire xformtmp108;
	assign xformtmp108 = ~xformtmp109;
	wire xformtmp272;
	assign xformtmp272 = xformtmp271 & xformtmp108;
	wire xformtmp269;
	assign xformtmp269 = ~xformtmp272;
	wire xformtmp275;
	assign xformtmp275 = xformtmp265 & xformtmp269;
	wire xformtmp232;
	assign xformtmp232 = in[28] & xformtmp218;
	wire xformtmp231;
	assign xformtmp231 = ~xformtmp232;
	wire xformtmp262;
	assign xformtmp262 = in[25] & xformtmp231;
	wire xformtmp187;
	assign xformtmp187 = in[26] & xformtmp164;
	wire xformtmp186;
	assign xformtmp186 = ~xformtmp187;
	wire xformtmp263;
	assign xformtmp263 = xformtmp262 & xformtmp186;
	wire xformtmp105;
	assign xformtmp105 = in[23] & xformtmp82;
	wire xformtmp104;
	assign xformtmp104 = ~xformtmp105;
	wire xformtmp264;
	assign xformtmp264 = xformtmp263 & xformtmp104;
	wire xformtmp261;
	assign xformtmp261 = ~xformtmp264;
	wire xformtmp276;
	assign xformtmp276 = xformtmp275 & xformtmp261;
	wire xformtmp230;
	assign xformtmp230 = in[24] & xformtmp218;
	wire xformtmp229;
	assign xformtmp229 = ~xformtmp230;
	wire xformtmp258;
	assign xformtmp258 = in[21] & xformtmp229;
	wire xformtmp185;
	assign xformtmp185 = in[22] & xformtmp164;
	wire xformtmp184;
	assign xformtmp184 = ~xformtmp185;
	wire xformtmp259;
	assign xformtmp259 = xformtmp258 & xformtmp184;
	wire xformtmp103;
	assign xformtmp103 = in[19] & xformtmp82;
	wire xformtmp102;
	assign xformtmp102 = ~xformtmp103;
	wire xformtmp260;
	assign xformtmp260 = xformtmp259 & xformtmp102;
	wire xformtmp257;
	assign xformtmp257 = ~xformtmp260;
	wire xformtmp277;
	assign xformtmp277 = xformtmp276 & xformtmp257;
	wire xformtmp228;
	assign xformtmp228 = in[20] & xformtmp218;
	wire xformtmp227;
	assign xformtmp227 = ~xformtmp228;
	wire xformtmp254;
	assign xformtmp254 = in[17] & xformtmp227;
	wire xformtmp182;
	assign xformtmp182 = in[18] & xformtmp164;
	wire xformtmp181;
	assign xformtmp181 = ~xformtmp182;
	wire xformtmp255;
	assign xformtmp255 = xformtmp254 & xformtmp181;
	wire xformtmp101;
	assign xformtmp101 = in[15] & xformtmp82;
	wire xformtmp100;
	assign xformtmp100 = ~xformtmp101;
	wire xformtmp256;
	assign xformtmp256 = xformtmp255 & xformtmp100;
	wire xformtmp253;
	assign xformtmp253 = ~xformtmp256;
	wire xformtmp278;
	assign xformtmp278 = xformtmp277 & xformtmp253;
	wire xformtmp226;
	assign xformtmp226 = in[16] & xformtmp218;
	wire xformtmp225;
	assign xformtmp225 = ~xformtmp226;
	wire xformtmp250;
	assign xformtmp250 = in[13] & xformtmp225;
	wire xformtmp179;
	assign xformtmp179 = in[14] & xformtmp164;
	wire xformtmp178;
	assign xformtmp178 = ~xformtmp179;
	wire xformtmp251;
	assign xformtmp251 = xformtmp250 & xformtmp178;
	wire xformtmp99;
	assign xformtmp99 = in[11] & xformtmp82;
	wire xformtmp98;
	assign xformtmp98 = ~xformtmp99;
	wire xformtmp252;
	assign xformtmp252 = xformtmp251 & xformtmp98;
	wire xformtmp249;
	assign xformtmp249 = ~xformtmp252;
	wire xformtmp279;
	assign xformtmp279 = xformtmp278 & xformtmp249;
	wire xformtmp224;
	assign xformtmp224 = in[12] & xformtmp218;
	wire xformtmp223;
	assign xformtmp223 = ~xformtmp224;
	wire xformtmp246;
	assign xformtmp246 = in[9] & xformtmp223;
	wire xformtmp176;
	assign xformtmp176 = in[10] & xformtmp164;
	wire xformtmp175;
	assign xformtmp175 = ~xformtmp176;
	wire xformtmp247;
	assign xformtmp247 = xformtmp246 & xformtmp175;
	wire xformtmp96;
	assign xformtmp96 = in[7] & xformtmp82;
	wire xformtmp95;
	assign xformtmp95 = ~xformtmp96;
	wire xformtmp248;
	assign xformtmp248 = xformtmp247 & xformtmp95;
	wire xformtmp245;
	assign xformtmp245 = ~xformtmp248;
	wire xformtmp280;
	assign xformtmp280 = xformtmp279 & xformtmp245;
	wire xformtmp222;
	assign xformtmp222 = in[8] & xformtmp218;
	wire xformtmp221;
	assign xformtmp221 = ~xformtmp222;
	wire xformtmp242;
	assign xformtmp242 = in[5] & xformtmp221;
	wire xformtmp173;
	assign xformtmp173 = in[6] & xformtmp164;
	wire xformtmp172;
	assign xformtmp172 = ~xformtmp173;
	wire xformtmp243;
	assign xformtmp243 = xformtmp242 & xformtmp172;
	wire xformtmp93;
	assign xformtmp93 = in[3] & xformtmp82;
	wire xformtmp92;
	assign xformtmp92 = ~xformtmp93;
	wire xformtmp244;
	assign xformtmp244 = xformtmp243 & xformtmp92;
	wire xformtmp241;
	assign xformtmp241 = ~xformtmp244;
	wire xformtmp274;
	assign xformtmp274 = xformtmp280 & xformtmp241;
	wire xformtmp285;
	assign xformtmp285 = xformtmp240 | xformtmp274;
	assign out[3] = ~xformtmp285;
	wire xformtmp287;
	assign xformtmp287 = xformtmp245 & xformtmp252;
	wire xformtmp286;
	assign xformtmp286 = ~xformtmp287;
	wire xformtmp299;
	assign xformtmp299 = xformtmp286 & xformtmp253;
	wire xformtmp300;
	assign xformtmp300 = xformtmp299 & xformtmp245;
	wire xformtmp301;
	assign xformtmp301 = xformtmp300 & xformtmp241;
	assign out[4] = ~xformtmp301;
	wire xformtmp289;
	assign xformtmp289 = xformtmp260 & xformtmp253;
	wire xformtmp290;
	assign xformtmp290 = xformtmp289 & xformtmp249;
	wire xformtmp291;
	assign xformtmp291 = xformtmp290 & xformtmp245;
	wire xformtmp288;
	assign xformtmp288 = ~xformtmp291;
	wire xformtmp293;
	assign xformtmp293 = xformtmp249 & xformtmp264;
	wire xformtmp294;
	assign xformtmp294 = xformtmp293 & xformtmp253;
	wire xformtmp292;
	assign xformtmp292 = ~xformtmp294;
	wire xformtmp302;
	assign xformtmp302 = xformtmp288 & xformtmp292;
	wire xformtmp303;
	assign xformtmp303 = xformtmp302 & xformtmp245;
	wire xformtmp304;
	assign xformtmp304 = xformtmp303 & xformtmp241;
	assign out[5] = ~xformtmp304;
	wire xformtmp296;
	assign xformtmp296 = xformtmp261 & xformtmp268;
	wire xformtmp297;
	assign xformtmp297 = xformtmp296 & xformtmp249;
	wire xformtmp298;
	assign xformtmp298 = xformtmp297 & xformtmp245;
	wire xformtmp295;
	assign xformtmp295 = ~xformtmp298;
	wire xformtmp305;
	assign xformtmp305 = xformtmp288 & xformtmp295;
	wire xformtmp306;
	assign xformtmp306 = xformtmp305 & xformtmp286;
	wire xformtmp307;
	assign xformtmp307 = xformtmp306 & xformtmp241;
	assign out[6] = ~xformtmp307;
endmodule

module tb();
    reg[6:0] results[1];
    reg[35:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%36b]", data[0]);
        #1
        $display("results = [%7b]", results[0]);
        $writememb("results.txt", results);
    end
endmodule

