module dut (out, in);
	output[79:0] out;
	input[149:0] in;
	wire origtmp1;
	wire origtmp2;
	wire origtmp3;
	wire origtmp4;
	wire origtmp5;
	wire origtmp6;
	wire origtmp7;
	wire origtmp8;
	wire origtmp9;
	wire origtmp10;
	wire origtmp11;
	wire origtmp12;
	wire origtmp13;
	wire origtmp14;
	wire origtmp15;
	wire origtmp16;
	wire origtmp17;
	wire origtmp18;
	wire origtmp19;
	wire origtmp20;
	wire origtmp21;
	wire origtmp22;
	wire origtmp23;
	wire origtmp24;
	wire origtmp25;
	wire origtmp26;
	wire origtmp27;
	wire origtmp28;
	wire origtmp29;
	wire origtmp30;
	wire origtmp31;
	wire origtmp32;
	wire origtmp33;
	wire origtmp34;
	wire origtmp35;
	wire origtmp36;
	wire origtmp37;
	wire origtmp38;
	wire origtmp39;
	wire origtmp40;
	wire origtmp41;
	wire origtmp42;
	wire origtmp43;
	wire origtmp44;
	wire origtmp45;
	wire origtmp46;
	wire origtmp47;
	wire origtmp48;
	wire origtmp49;
	wire origtmp50;
	wire origtmp51;
	wire origtmp52;
	wire origtmp53;
	wire origtmp54;
	wire origtmp55;
	wire origtmp56;
	wire origtmp57;
	wire origtmp58;
	wire origtmp59;
	wire origtmp60;
	wire origtmp61;
	wire origtmp62;
	wire origtmp63;
	wire origtmp64;
	wire origtmp65;
	wire origtmp66;
	wire origtmp67;
	wire origtmp68;
	wire origtmp69;
	wire origtmp70;
	wire origtmp71;
	wire origtmp72;
	wire origtmp73;
	wire origtmp74;
	wire origtmp75;
	wire origtmp76;
	wire origtmp77;
	wire origtmp78;
	wire origtmp79;
	wire origtmp80;
	wire origtmp81;
	wire origtmp82;
	wire origtmp83;
	wire origtmp84;
	wire origtmp85;
	wire origtmp86;
	wire origtmp87;
	wire origtmp88;
	wire origtmp89;
	wire origtmp90;
	wire origtmp91;
	wire origtmp92;
	wire origtmp93;
	wire origtmp94;
	wire origtmp95;
	wire origtmp96;
	wire origtmp97;
	wire origtmp98;
	wire origtmp99;
	wire origtmp100;
	wire origtmp101;
	wire origtmp102;
	wire origtmp103;
	wire origtmp104;
	wire origtmp105;
	wire origtmp106;
	wire origtmp107;
	wire origtmp108;
	wire origtmp109;
	wire origtmp110;
	wire origtmp111;
	wire origtmp112;
	wire origtmp113;
	wire origtmp114;
	wire origtmp115;
	wire origtmp116;
	wire origtmp117;
	wire origtmp118;
	wire origtmp119;
	wire origtmp120;
	wire origtmp121;
	wire origtmp122;
	wire origtmp123;
	wire origtmp124;
	wire origtmp125;
	wire origtmp126;
	wire origtmp127;
	wire origtmp128;
	wire origtmp129;
	wire origtmp130;
	wire origtmp131;
	wire origtmp132;
	wire origtmp133;
	wire origtmp134;
	wire origtmp135;
	wire origtmp136;
	wire origtmp137;
	wire origtmp138;
	wire origtmp139;
	wire origtmp140;
	wire origtmp141;
	wire origtmp142;
	wire origtmp143;
	wire origtmp144;
	wire origtmp145;
	wire origtmp146;
	wire origtmp147;
	wire origtmp148;
	wire origtmp149;
	wire origtmp150;
	wire origtmp151;
	wire origtmp152;
	wire origtmp153;
	wire origtmp154;
	wire origtmp155;
	wire origtmp156;
	wire origtmp157;
	wire origtmp158;
	wire origtmp159;
	wire origtmp160;
	wire origtmp161;
	wire origtmp162;
	wire origtmp163;
	wire origtmp164;
	wire origtmp165;
	wire origtmp166;
	wire origtmp167;
	wire origtmp168;
	wire origtmp169;
	wire origtmp170;
	wire origtmp171;
	wire origtmp172;
	wire origtmp173;
	wire origtmp174;
	wire origtmp175;
	wire origtmp176;
	wire origtmp177;
	wire origtmp178;
	wire origtmp179;
	wire origtmp180;
	wire origtmp181;
	wire origtmp182;
	wire origtmp183;
	wire origtmp184;
	wire origtmp185;
	wire origtmp186;
	wire origtmp187;
	wire origtmp188;
	wire origtmp189;
	wire origtmp190;
	wire origtmp191;
	wire origtmp192;
	wire origtmp193;
	wire origtmp194;
	wire origtmp195;
	wire origtmp196;
	wire origtmp197;
	wire origtmp198;
	wire origtmp199;
	wire origtmp200;
	wire origtmp201;
	wire origtmp202;
	wire origtmp203;
	wire origtmp204;
	wire origtmp205;
	wire origtmp206;
	wire origtmp207;
	wire origtmp208;
	wire origtmp209;
	wire origtmp210;
	wire origtmp211;
	wire origtmp212;
	wire origtmp213;
	wire origtmp214;
	wire origtmp215;
	wire origtmp216;
	wire origtmp217;
	wire origtmp218;
	wire origtmp219;
	wire origtmp220;
	wire origtmp221;
	assign origtmp207 = 1'b1;
	assign out[61] = origtmp209 & 1'b1;
	assign origtmp191 = 1'b1;
	assign out[60] = 1'b0;
	assign origtmp44 = in[116] | in[115];
	assign origtmp210 = 1'b0;
	assign origtmp68 = 1'b0 ^ origtmp108;
	assign out[79] = origtmp221 ^ 1'b0;
	assign origtmp189 = 1'b0 | 1'b0;
	assign origtmp112 = in[108] & in[113];
	assign origtmp53 = ~in[83];
	assign origtmp60 = ~in[145];
	assign origtmp107 = in[27] ^ origtmp65;
	assign out[67] = 1'b0 & 1'b0;
	assign out[12] = origtmp181 | origtmp181;
	assign out[57] = 1'b1;
	assign origtmp63 = origtmp85 ^ origtmp101;
	assign out[66] = origtmp214 & origtmp214;
	assign origtmp168 = in[60] & in[34];
	assign origtmp172 = 1'b0 & origtmp173;
	assign origtmp159 = in[0] & in[94];
	assign origtmp178 = in[22] | in[54];
	assign out[10] = origtmp180;
	assign origtmp47 = origtmp37 & in[2];
	assign origtmp208 = 1'b0 | 1'b1;
	assign origtmp169 = origtmp139 | origtmp129;
	assign origtmp188 = 1'b0;
	assign origtmp91 = in[87] & in[18];
	assign out[68] = 1'b1;
	assign origtmp138 = in[131] ^ in[77];
	assign origtmp114 = origtmp123 | origtmp76;
	assign origtmp119 = origtmp106 & in[110];
	assign origtmp174 = in[70] ^ origtmp177;
	assign origtmp31 = in[142] & in[20];
	assign out[63] = origtmp211 | origtmp211;
	assign origtmp94 = in[15] | origtmp96;
	assign out[55] = origtmp207 ^ 1'b1;
	assign origtmp220 = 1'b1 | 1'b1;
	assign origtmp136 = in[57] | in[9];
	assign out[49] = origtmp204 & 1'b0;
	assign origtmp80 = in[103] & in[87];
	assign origtmp105 = in[40] | in[11];
	assign origtmp11 = origtmp47 | origtmp15;
	assign origtmp55 = origtmp49 & origtmp29;
	assign origtmp59 = origtmp75 ^ origtmp97;
	assign out[56] = 1'b0 | 1'b0;
	assign origtmp147 = in[50] ^ in[8];
	assign origtmp153 = in[129] & in[14];
	assign out[78] = ~origtmp220;
	assign origtmp142 = origtmp146 | origtmp141;
	assign origtmp64 = in[52] | in[136];
	assign origtmp66 = origtmp74 | origtmp79;
	assign origtmp32 = in[71] | in[138];
	assign origtmp201 = 1'b0 & 1'b0;
	assign origtmp139 = origtmp170 & origtmp145;
	assign out[59] = 1'b1 ^ origtmp208;
	assign origtmp158 = origtmp161 & in[95];
	assign origtmp148 = origtmp143 | origtmp153;
	assign origtmp152 = origtmp148 ^ origtmp155;
	assign origtmp127 = in[120] | in[13];
	assign origtmp56 = origtmp59 | origtmp104;
	assign origtmp109 = in[63] | in[45];
	assign out[5] = origtmp174 ^ origtmp176;
	assign origtmp40 = in[142] ^ in[62];
	assign origtmp111 = in[61] | in[81];
	assign out[23] = origtmp188;
	assign origtmp205 = ~1'b1;
	assign origtmp16 = origtmp2 ^ origtmp1;
	assign origtmp96 = in[25] ^ in[61];
	assign origtmp102 = origtmp119 | origtmp88;
	assign origtmp89 = origtmp66 ^ origtmp112;
	assign origtmp177 = in[66] | origtmp175;
	assign out[74] = 1'b1;
	assign origtmp171 = origtmp166 & origtmp131;
	assign origtmp196 = 1'b1;
	assign origtmp28 = in[26] | in[137];
	assign origtmp14 = in[124] & in[121];
	assign origtmp38 = in[119] & in[107];
	assign origtmp15 = origtmp24 | origtmp20;
	assign origtmp135 = origtmp162 & in[75];
	assign origtmp209 = 1'b1 ^ 1'b0;
	assign out[62] = origtmp210;
	assign origtmp71 = in[18] & in[113];
	assign origtmp176 = in[66] & in[147];
	assign out[65] = origtmp213 | origtmp213;
	assign origtmp12 = in[79] | origtmp7;
	assign out[42] = origtmp199;
	assign origtmp128 = origtmp167 | origtmp159;
	assign out[39] = origtmp197 ^ origtmp197;
	assign origtmp87 = origtmp84 & origtmp56;
	assign out[24] = 1'b1;
	assign origtmp57 = origtmp77 ^ origtmp82;
	assign origtmp9 = origtmp44 ^ origtmp32;
	assign origtmp211 = ~1'b0;
	assign origtmp104 = in[143] | origtmp121;
	assign out[19] = ~origtmp186;
	assign out[58] = 1'b0 | 1'b1;
	assign origtmp150 = in[104] & origtmp140;
	assign out[27] = origtmp190 ^ origtmp190;
	assign out[64] = origtmp212 & origtmp212;
	assign origtmp212 = 1'b0;
	assign origtmp50 = origtmp22 & origtmp8;
	assign origtmp95 = origtmp87 | origtmp118;
	assign origtmp115 = in[46] & origtmp100;
	assign origtmp145 = in[146] & origtmp142;
	assign origtmp170 = in[23] | origtmp168;
	assign out[9] = 1'b1;
	assign out[50] = origtmp205 & origtmp205;
	assign out[26] = 1'b1 ^ 1'b1;
	assign origtmp156 = in[139] | in[111];
	assign origtmp213 = ~1'b0;
	assign origtmp10 = in[19] | in[24];
	assign origtmp110 = in[55] ^ in[15];
	assign origtmp22 = origtmp52 | in[47];
	assign origtmp43 = origtmp33 ^ origtmp18;
	assign origtmp195 = 1'b1 ^ 1'b0;
	assign out[31] = origtmp193 ^ origtmp193;
	assign origtmp106 = origtmp113 | in[97];
	assign out[28] = origtmp191 | origtmp191;
	assign origtmp37 = in[78] & in[53];
	assign out[4] = origtmp172 & in[21];
	assign origtmp131 = in[5] & origtmp169;
	assign origtmp13 = origtmp35 ^ in[24];
	assign origtmp103 = origtmp73 ^ origtmp95;
	assign origtmp23 = origtmp25 | in[62];
	assign out[47] = ~1'b1;
	assign out[40] = 1'b1 & origtmp198;
	assign origtmp126 = in[109] & in[144];
	assign origtmp84 = in[113] & 1'b1;
	assign out[70] = origtmp216 ^ origtmp216;
	assign origtmp39 = origtmp10 | origtmp13;
	assign origtmp21 = origtmp39 ^ origtmp48;
	assign out[53] = 1'b1 & 1'b0;
	assign out[54] = 1'b0 ^ 1'b1;
	assign origtmp90 = origtmp58 ^ origtmp105;
	assign origtmp183 = 1'b1 | 1'b1;
	assign origtmp100 = in[7] ^ in[29];
	assign origtmp26 = origtmp30 & origtmp46;
	assign origtmp86 = in[93] & origtmp111;
	assign out[11] = 1'b0 | 1'b1;
	assign origtmp73 = in[69] | in[68];
	assign out[69] = 1'b1 & origtmp215;
	assign out[25] = ~origtmp189;
	assign origtmp143 = origtmp163 ^ in[16];
	assign origtmp101 = origtmp61 & origtmp72;
	assign origtmp190 = ~1'b0;
	assign origtmp20 = origtmp27 & in[91];
	assign out[71] = origtmp217 ^ 1'b0;
	assign out[3] = origtmp134 | origtmp144;
	assign origtmp166 = in[86] ^ origtmp150;
	assign origtmp155 = origtmp157 ^ origtmp133;
	assign origtmp3 = in[128] & origtmp26;
	assign out[21] = 1'b0 ^ 1'b0;
	assign origtmp161 = origtmp128 & in[48];
	assign origtmp92 = in[41] | in[45];
	assign origtmp124 = origtmp102 | in[45];
	assign out[14] = 1'b0 | origtmp183;
	assign origtmp48 = in[142] & in[123];
	assign out[34] = origtmp195 & 1'b1;
	assign origtmp121 = origtmp107 ^ in[25];
	assign out[51] = 1'b1;
	assign out[75] = 1'b0 & origtmp219;
	assign origtmp187 = 1'b0;
	assign origtmp137 = origtmp171 ^ origtmp138;
	assign origtmp78 = in[143] & origtmp92;
	assign origtmp67 = in[45] & in[101];
	assign origtmp160 = in[73] | in[95];
	assign origtmp52 = in[39] ^ in[124];
	assign origtmp144 = origtmp132 & origtmp154;
	assign out[72] = ~1'b0;
	assign origtmp118 = origtmp60 | origtmp117;
	assign out[30] = origtmp192 ^ 1'b0;
	assign out[76] = 1'b1;
	assign origtmp186 = ~1'b1;
	assign out[1] = origtmp63 | origtmp103;
	assign origtmp193 = ~1'b1;
	assign origtmp29 = origtmp34 ^ origtmp42;
	assign origtmp62 = origtmp110 ^ in[112];
	assign origtmp216 = ~1'b0;
	assign origtmp184 = 1'b1 & 1'b1;
	assign origtmp146 = origtmp135 | in[106];
	assign origtmp203 = 1'b0 & 1'b1;
	assign origtmp6 = in[85] ^ origtmp5;
	assign origtmp36 = in[72] & origtmp41;
	assign origtmp162 = in[28] | in[102];
	assign out[18] = origtmp185 ^ 1'b0;
	assign out[16] = 1'b0;
	assign origtmp4 = in[64] & in[96];
	assign origtmp221 = in[100] | in[100];
	assign origtmp77 = in[133] & in[136];
	assign out[41] = ~1'b1;
	assign out[46] = 1'b0;
	assign origtmp141 = in[89] | in[135];
	assign origtmp54 = origtmp4 & in[31];
	assign origtmp19 = in[82] & in[30];
	assign origtmp1 = origtmp28 & origtmp53;
	assign origtmp173 = in[134] | in[49];
	assign origtmp125 = origtmp127 ^ origtmp126;
	assign origtmp7 = in[107] & in[17];
	assign origtmp133 = origtmp164 | in[4];
	assign origtmp219 = 1'b0;
	assign out[36] = 1'b0 & 1'b1;
	assign origtmp132 = origtmp158 & origtmp165;
	assign origtmp198 = 1'b1 & 1'b0;
	assign origtmp181 = 1'b0;
	assign origtmp167 = in[99] ^ in[67];
	assign origtmp82 = origtmp86 & origtmp83;
	assign origtmp214 = 1'b0 & 1'b1;
	assign origtmp69 = in[40] & in[46];
	assign origtmp157 = origtmp130 | in[8];
	assign origtmp74 = in[130] & origtmp71;
	assign origtmp72 = origtmp120 | origtmp64;
	assign out[13] = origtmp182;
	assign origtmp30 = origtmp40 | in[141];
	assign origtmp97 = origtmp62 & in[15];
	assign origtmp99 = origtmp98 & in[10];
	assign out[33] = 1'b0 ^ origtmp194;
	assign out[20] = 1'b0 | 1'b1;
	assign out[15] = 1'b0 & 1'b1;
	assign origtmp194 = 1'b1 & 1'b0;
	assign origtmp130 = in[56] | in[105];
	assign origtmp192 = 1'b0;
	assign out[22] = origtmp187;
	assign out[48] = origtmp203 & origtmp203;
	assign origtmp17 = origtmp16 ^ origtmp21;
	assign origtmp182 = 1'b1;
	assign origtmp25 = in[12] ^ in[71];
	assign origtmp197 = 1'b0 & 1'b0;
	assign origtmp83 = origtmp99 & in[143];
	assign origtmp88 = origtmp91 & origtmp109;
	assign origtmp27 = origtmp9 & origtmp6;
	assign origtmp199 = 1'b1;
	assign origtmp2 = origtmp19 & in[35];
	assign origtmp165 = in[38] | origtmp160;
	assign origtmp204 = 1'b0 ^ 1'b0;
	assign out[45] = origtmp202 & 1'b1;
	assign out[43] = ~origtmp200;
	assign origtmp33 = in[64] ^ origtmp14;
	assign origtmp5 = origtmp38 ^ in[35];
	assign origtmp79 = in[15] | origtmp122;
	assign origtmp116 = in[27] & in[45];
	assign origtmp215 = 1'b1 | 1'b1;
	assign out[37] = 1'b1;
	assign origtmp140 = in[132] ^ in[37];
	assign origtmp206 = 1'b0;
	assign origtmp70 = origtmp89 & origtmp67;
	assign out[52] = 1'b0 & origtmp206;
	assign origtmp24 = origtmp31 | origtmp23;
	assign origtmp49 = origtmp50 & origtmp36;
	assign origtmp45 = origtmp17 | origtmp55;
	assign origtmp18 = in[6] ^ in[91];
	assign origtmp34 = in[33] | in[32];
	assign origtmp46 = origtmp11 | origtmp51;
	assign out[8] = 1'b0;
	assign origtmp81 = origtmp93 & origtmp70;
	assign origtmp42 = origtmp54 ^ in[149];
	assign origtmp75 = in[148] ^ origtmp80;
	assign origtmp164 = origtmp151 | origtmp156;
	assign origtmp154 = origtmp147 & origtmp149;
	assign origtmp65 = in[114] ^ in[127];
	assign origtmp58 = in[114] ^ origtmp116;
	assign origtmp8 = in[43] | in[76];
	assign origtmp180 = 1'b0;
	assign out[35] = 1'b0;
	assign origtmp179 = 1'b0;
	assign origtmp98 = ~in[90];
	assign origtmp123 = origtmp69 ^ in[58];
	assign origtmp108 = in[125] | in[88];
	assign origtmp200 = 1'b0 & 1'b1;
	assign origtmp134 = origtmp152 ^ origtmp137;
	assign out[77] = 1'b1 ^ 1'b0;
	assign origtmp202 = 1'b1;
	assign origtmp93 = origtmp57 & origtmp115;
	assign origtmp85 = origtmp124 | origtmp94;
	assign out[0] = origtmp45 & origtmp3;
	assign origtmp129 = origtmp136 ^ in[65];
	assign origtmp217 = ~1'b0;
	assign origtmp175 = in[118] & in[66];
	assign origtmp163 = in[42] | in[80];
	assign origtmp122 = in[3] | in[29];
	assign origtmp151 = in[126] & in[36];
	assign origtmp149 = in[92] & in[98];
	assign out[32] = 1'b0;
	assign out[38] = origtmp196 & 1'b0;
	assign origtmp51 = origtmp43 & in[140];
	assign origtmp117 = origtmp78 | in[113];
	assign out[17] = origtmp184 | origtmp184;
	assign out[29] = 1'b1 ^ 1'b0;
	assign origtmp41 = origtmp12 | in[117];
	assign origtmp218 = 1'b0;
	assign origtmp185 = 1'b1 & 1'b1;
	assign origtmp120 = origtmp90 & origtmp68;
	assign origtmp35 = in[122] & in[1];
	assign out[73] = origtmp218 & origtmp218;
	assign out[2] = in[51] & origtmp125;
	assign out[7] = origtmp179;
	assign out[6] = origtmp178 | in[84];
	assign out[44] = origtmp201 ^ origtmp201;
	assign origtmp76 = in[59] | in[108];
	assign origtmp61 = origtmp81 | origtmp114;
	assign origtmp113 = in[44] | in[74];
endmodule

module tb();
    reg[79:0] results[1];
    reg[149:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%150b]", data[0]);
        #1
        $display("results = [%80b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
