module dut (out, in);
	output[1:0] out;
	input[1:0] in;
	wire origtmp1;
	wire origtmp2;
	wire origtmp3;
	wire origtmp4;
	wire origtmp5;
	wire origtmp6;
	wire origtmp7;
	wire origtmp8;
	wire origtmp9;
	wire origtmp10;
	wire origtmp11;
	wire origtmp12;
	wire origtmp13;
	wire origtmp14;
	wire origtmp15;
	wire origtmp16;
	wire origtmp17;
	wire origtmp18;
	wire origtmp19;
	wire origtmp20;
	wire origtmp21;
	wire origtmp22;
	wire origtmp23;
	wire origtmp24;
	wire origtmp25;
	wire origtmp26;
	wire origtmp27;
	wire origtmp28;
	wire origtmp29;
	wire origtmp30;
	wire origtmp31;
	wire origtmp32;
	wire origtmp33;
	wire origtmp34;
	wire origtmp35;
	wire origtmp36;
	wire origtmp37;
	wire origtmp38;
	wire origtmp39;
	wire origtmp40;
	wire origtmp41;
	wire origtmp42;
	wire origtmp43;
	wire origtmp44;
	wire origtmp45;
	wire origtmp46;
	wire origtmp47;
	wire origtmp48;
	wire origtmp49;
	wire origtmp50;
	assign origtmp1 = ~in[0];
	assign origtmp2 = origtmp1;
	assign origtmp3 = origtmp2 ^ 1'b0;
	assign origtmp4 = origtmp3 | 1'b0;
	assign origtmp5 = origtmp4 & 1'b1;
	assign origtmp6 = origtmp5 ^ 1'b0;
	assign origtmp7 = origtmp6 ^ 1'b1;
	assign origtmp8 = origtmp7 ^ 1'b1;
	assign origtmp9 = origtmp8 | 1'b0;
	assign origtmp10 = origtmp9 ^ 1'b0;
	assign origtmp11 = origtmp10 ^ 1'b0;
	assign origtmp12 = origtmp11 ^ 1'b1;
	assign origtmp13 = origtmp12 | 1'b0;
	assign origtmp14 = origtmp13;
	assign origtmp15 = ~origtmp14;
	assign origtmp16 = origtmp15 ^ 1'b1;
	assign origtmp17 = origtmp16 & 1'b1;
	assign origtmp18 = origtmp17 ^ 1'b1;
	assign origtmp19 = origtmp18 ^ 1'b0;
	assign origtmp20 = origtmp19 | 1'b0;
	assign origtmp21 = origtmp20;
	assign origtmp22 = origtmp21;
	assign origtmp23 = origtmp22;
	assign origtmp24 = ~origtmp23;
	assign origtmp25 = origtmp24 | 1'b0;
	assign origtmp26 = origtmp25 | 1'b0;
	assign origtmp27 = ~origtmp26;
	assign origtmp28 = origtmp27;
	assign origtmp29 = origtmp28 ^ 1'b0;
	assign origtmp30 = ~origtmp29;
	assign origtmp31 = origtmp30 & 1'b1;
	assign origtmp32 = origtmp31 ^ 1'b0;
	assign origtmp33 = origtmp32 ^ 1'b1;
	assign origtmp34 = origtmp33 & 1'b1;
	assign origtmp35 = origtmp34 | 1'b0;
	assign origtmp36 = origtmp35;
	assign origtmp37 = origtmp36 ^ 1'b0;
	assign origtmp38 = ~origtmp37;
	assign origtmp39 = origtmp38 & 1'b1;
	assign origtmp40 = origtmp39 ^ 1'b1;
	assign origtmp41 = origtmp40 ^ 1'b0;
	assign origtmp42 = ~origtmp41;
	assign origtmp43 = origtmp42 ^ 1'b1;
	assign origtmp44 = origtmp43;
	assign origtmp45 = origtmp44 & 1'b1;
	assign origtmp46 = origtmp45 & 1'b1;
	assign origtmp47 = origtmp46 ^ 1'b0;
	assign origtmp48 = ~origtmp47;
	assign origtmp49 = origtmp48 ^ 1'b1;
	assign origtmp50 = origtmp49 ^ 1'b0;
	assign out[0] = origtmp50 ^ 1'b0;
	assign out[1] = origtmp50 ^ in[1];
endmodule

module tb();
    reg[1:0] results[1];
    reg[1:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%2b]", data[0]);
        #1
        $display("results = [%2b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
