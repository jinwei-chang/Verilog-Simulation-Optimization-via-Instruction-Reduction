module dut (out, in);
	output[79:0] out;
	input[149:0] in;
	wire xformtmp19;
	assign xformtmp19 = in[82] & in[30];
	wire xformtmp2;
	assign xformtmp2 = xformtmp19 & in[35];
	wire xformtmp28;
	assign xformtmp28 = in[26] | in[137];
	wire xformtmp53;
	assign xformtmp53 = ~in[83];
	wire xformtmp1;
	assign xformtmp1 = xformtmp28 & xformtmp53;
	wire xformtmp16;
	assign xformtmp16 = xformtmp2 ^ xformtmp1;
	wire xformtmp10;
	assign xformtmp10 = in[19] | in[24];
	wire xformtmp35;
	assign xformtmp35 = in[122] & in[1];
	wire xformtmp13;
	assign xformtmp13 = xformtmp35 ^ in[24];
	wire xformtmp39;
	assign xformtmp39 = xformtmp10 | xformtmp13;
	wire xformtmp48;
	assign xformtmp48 = in[142] & in[123];
	wire xformtmp21;
	assign xformtmp21 = xformtmp39 ^ xformtmp48;
	wire xformtmp17;
	assign xformtmp17 = xformtmp16 ^ xformtmp21;
	wire xformtmp52;
	assign xformtmp52 = in[39] ^ in[124];
	wire xformtmp22;
	assign xformtmp22 = xformtmp52 | in[47];
	wire xformtmp8;
	assign xformtmp8 = in[43] | in[76];
	wire xformtmp50;
	assign xformtmp50 = xformtmp22 & xformtmp8;
	wire xformtmp7;
	assign xformtmp7 = in[107] & in[17];
	wire xformtmp12;
	assign xformtmp12 = in[79] | xformtmp7;
	wire xformtmp41;
	assign xformtmp41 = xformtmp12 | in[117];
	wire xformtmp36;
	assign xformtmp36 = in[72] & xformtmp41;
	wire xformtmp49;
	assign xformtmp49 = xformtmp50 & xformtmp36;
	wire xformtmp34;
	assign xformtmp34 = in[33] | in[32];
	wire xformtmp4;
	assign xformtmp4 = in[64] & in[96];
	wire xformtmp54;
	assign xformtmp54 = xformtmp4 & in[31];
	wire xformtmp42;
	assign xformtmp42 = xformtmp54 ^ in[149];
	wire xformtmp29;
	assign xformtmp29 = xformtmp34 ^ xformtmp42;
	wire xformtmp55;
	assign xformtmp55 = xformtmp49 & xformtmp29;
	wire xformtmp45;
	assign xformtmp45 = xformtmp17 | xformtmp55;
	wire xformtmp40;
	assign xformtmp40 = in[142] ^ in[62];
	wire xformtmp30;
	assign xformtmp30 = xformtmp40 | in[141];
	wire xformtmp37;
	assign xformtmp37 = in[78] & in[53];
	wire xformtmp47;
	assign xformtmp47 = xformtmp37 & in[2];
	wire xformtmp31;
	assign xformtmp31 = in[142] & in[20];
	wire xformtmp25;
	assign xformtmp25 = in[12] ^ in[71];
	wire xformtmp23;
	assign xformtmp23 = xformtmp25 | in[62];
	wire xformtmp24;
	assign xformtmp24 = xformtmp31 | xformtmp23;
	wire xformtmp44;
	assign xformtmp44 = in[116] | in[115];
	wire xformtmp32;
	assign xformtmp32 = in[71] | in[138];
	wire xformtmp9;
	assign xformtmp9 = xformtmp44 ^ xformtmp32;
	wire xformtmp38;
	assign xformtmp38 = in[119] & in[107];
	wire xformtmp5;
	assign xformtmp5 = xformtmp38 ^ in[35];
	wire xformtmp6;
	assign xformtmp6 = in[85] ^ xformtmp5;
	wire xformtmp27;
	assign xformtmp27 = xformtmp9 & xformtmp6;
	wire xformtmp20;
	assign xformtmp20 = xformtmp27 & in[91];
	wire xformtmp15;
	assign xformtmp15 = xformtmp24 | xformtmp20;
	wire xformtmp11;
	assign xformtmp11 = xformtmp47 | xformtmp15;
	wire xformtmp14;
	assign xformtmp14 = in[124] & in[121];
	wire xformtmp33;
	assign xformtmp33 = in[64] ^ xformtmp14;
	wire xformtmp18;
	assign xformtmp18 = in[6] ^ in[91];
	wire xformtmp43;
	assign xformtmp43 = xformtmp33 ^ xformtmp18;
	wire xformtmp51;
	assign xformtmp51 = xformtmp43 & in[140];
	wire xformtmp46;
	assign xformtmp46 = xformtmp11 | xformtmp51;
	wire xformtmp26;
	assign xformtmp26 = xformtmp30 & xformtmp46;
	wire xformtmp3;
	assign xformtmp3 = in[128] & xformtmp26;
	assign out[0] = xformtmp45 & xformtmp3;
	wire xformtmp113;
	assign xformtmp113 = in[44] | in[74];
	wire xformtmp106;
	assign xformtmp106 = xformtmp113 | in[97];
	wire xformtmp119;
	assign xformtmp119 = xformtmp106 & in[110];
	wire xformtmp91;
	assign xformtmp91 = in[87] & in[18];
	wire xformtmp109;
	assign xformtmp109 = in[63] | in[45];
	wire xformtmp88;
	assign xformtmp88 = xformtmp91 & xformtmp109;
	wire xformtmp102;
	assign xformtmp102 = xformtmp119 | xformtmp88;
	wire xformtmp124;
	assign xformtmp124 = xformtmp102 | in[45];
	wire xformtmp96;
	assign xformtmp96 = in[25] ^ in[61];
	wire xformtmp94;
	assign xformtmp94 = in[15] | xformtmp96;
	wire xformtmp85;
	assign xformtmp85 = xformtmp124 | xformtmp94;
	wire xformtmp77;
	assign xformtmp77 = in[133] & in[136];
	wire xformtmp111;
	assign xformtmp111 = in[61] | in[81];
	wire xformtmp86;
	assign xformtmp86 = in[93] & xformtmp111;
	wire xformtmp98;
	assign xformtmp98 = ~in[90];
	wire xformtmp99;
	assign xformtmp99 = xformtmp98 & in[10];
	wire xformtmp83;
	assign xformtmp83 = xformtmp99 & in[143];
	wire xformtmp82;
	assign xformtmp82 = xformtmp86 & xformtmp83;
	wire xformtmp57;
	assign xformtmp57 = xformtmp77 ^ xformtmp82;
	wire xformtmp100;
	assign xformtmp100 = in[7] ^ in[29];
	wire xformtmp115;
	assign xformtmp115 = in[46] & xformtmp100;
	wire xformtmp93;
	assign xformtmp93 = xformtmp57 & xformtmp115;
	wire xformtmp71;
	assign xformtmp71 = in[18] & in[113];
	wire xformtmp74;
	assign xformtmp74 = in[130] & xformtmp71;
	wire xformtmp122;
	assign xformtmp122 = in[3] | in[29];
	wire xformtmp79;
	assign xformtmp79 = in[15] | xformtmp122;
	wire xformtmp66;
	assign xformtmp66 = xformtmp74 | xformtmp79;
	wire xformtmp112;
	assign xformtmp112 = in[108] & in[113];
	wire xformtmp89;
	assign xformtmp89 = xformtmp66 ^ xformtmp112;
	wire xformtmp67;
	assign xformtmp67 = in[45] & in[101];
	wire xformtmp70;
	assign xformtmp70 = xformtmp89 & xformtmp67;
	wire xformtmp81;
	assign xformtmp81 = xformtmp93 & xformtmp70;
	wire xformtmp69;
	assign xformtmp69 = in[40] & in[46];
	wire xformtmp123;
	assign xformtmp123 = xformtmp69 ^ in[58];
	wire xformtmp76;
	assign xformtmp76 = in[59] | in[108];
	wire xformtmp114;
	assign xformtmp114 = xformtmp123 | xformtmp76;
	wire xformtmp61;
	assign xformtmp61 = xformtmp81 | xformtmp114;
	wire xformtmp116;
	assign xformtmp116 = in[27] & in[45];
	wire xformtmp58;
	assign xformtmp58 = in[114] ^ xformtmp116;
	wire xformtmp105;
	assign xformtmp105 = in[40] | in[11];
	wire xformtmp90;
	assign xformtmp90 = xformtmp58 ^ xformtmp105;
	wire xformtmp108;
	assign xformtmp108 = in[125] | in[88];
	wire xformtmp120;
	assign xformtmp120 = xformtmp90 & xformtmp108;
	wire xformtmp64;
	assign xformtmp64 = in[52] | in[136];
	wire xformtmp72;
	assign xformtmp72 = xformtmp120 | xformtmp64;
	wire xformtmp101;
	assign xformtmp101 = xformtmp61 & xformtmp72;
	wire xformtmp63;
	assign xformtmp63 = xformtmp85 ^ xformtmp101;
	wire xformtmp73;
	assign xformtmp73 = in[69] | in[68];
	wire xformtmp80;
	assign xformtmp80 = in[103] & in[87];
	wire xformtmp75;
	assign xformtmp75 = in[148] ^ xformtmp80;
	wire xformtmp110;
	assign xformtmp110 = in[55] ^ in[15];
	wire xformtmp62;
	assign xformtmp62 = xformtmp110 ^ in[112];
	wire xformtmp97;
	assign xformtmp97 = xformtmp62 & in[15];
	wire xformtmp59;
	assign xformtmp59 = xformtmp75 ^ xformtmp97;
	wire xformtmp65;
	assign xformtmp65 = in[114] ^ in[127];
	wire xformtmp107;
	assign xformtmp107 = in[27] ^ xformtmp65;
	wire xformtmp121;
	assign xformtmp121 = xformtmp107 ^ in[25];
	wire xformtmp104;
	assign xformtmp104 = in[143] | xformtmp121;
	wire xformtmp56;
	assign xformtmp56 = xformtmp59 | xformtmp104;
	wire xformtmp87;
	assign xformtmp87 = in[113] & xformtmp56;
	wire xformtmp60;
	assign xformtmp60 = ~in[145];
	wire xformtmp92;
	assign xformtmp92 = in[41] | in[45];
	wire xformtmp78;
	assign xformtmp78 = in[143] & xformtmp92;
	wire xformtmp117;
	assign xformtmp117 = xformtmp78 | in[113];
	wire xformtmp118;
	assign xformtmp118 = xformtmp60 | xformtmp117;
	wire xformtmp95;
	assign xformtmp95 = xformtmp87 | xformtmp118;
	wire xformtmp103;
	assign xformtmp103 = xformtmp73 ^ xformtmp95;
	assign out[1] = xformtmp63 | xformtmp103;
	wire xformtmp127;
	assign xformtmp127 = in[120] | in[13];
	wire xformtmp126;
	assign xformtmp126 = in[109] & in[144];
	wire xformtmp125;
	assign xformtmp125 = xformtmp127 ^ xformtmp126;
	assign out[2] = in[51] & xformtmp125;
	wire xformtmp163;
	assign xformtmp163 = in[42] | in[80];
	wire xformtmp143;
	assign xformtmp143 = xformtmp163 ^ in[16];
	wire xformtmp153;
	assign xformtmp153 = in[129] & in[14];
	wire xformtmp148;
	assign xformtmp148 = xformtmp143 | xformtmp153;
	wire xformtmp130;
	assign xformtmp130 = in[56] | in[105];
	wire xformtmp157;
	assign xformtmp157 = xformtmp130 | in[8];
	wire xformtmp151;
	assign xformtmp151 = in[126] & in[36];
	wire xformtmp156;
	assign xformtmp156 = in[139] | in[111];
	wire xformtmp164;
	assign xformtmp164 = xformtmp151 | xformtmp156;
	wire xformtmp133;
	assign xformtmp133 = xformtmp164 | in[4];
	wire xformtmp155;
	assign xformtmp155 = xformtmp157 ^ xformtmp133;
	wire xformtmp152;
	assign xformtmp152 = xformtmp148 ^ xformtmp155;
	wire xformtmp140;
	assign xformtmp140 = in[132] ^ in[37];
	wire xformtmp150;
	assign xformtmp150 = in[104] & xformtmp140;
	wire xformtmp166;
	assign xformtmp166 = in[86] ^ xformtmp150;
	wire xformtmp168;
	assign xformtmp168 = in[60] & in[34];
	wire xformtmp170;
	assign xformtmp170 = in[23] | xformtmp168;
	wire xformtmp162;
	assign xformtmp162 = in[28] | in[102];
	wire xformtmp135;
	assign xformtmp135 = xformtmp162 & in[75];
	wire xformtmp146;
	assign xformtmp146 = xformtmp135 | in[106];
	wire xformtmp141;
	assign xformtmp141 = in[89] | in[135];
	wire xformtmp142;
	assign xformtmp142 = xformtmp146 | xformtmp141;
	wire xformtmp145;
	assign xformtmp145 = in[146] & xformtmp142;
	wire xformtmp139;
	assign xformtmp139 = xformtmp170 & xformtmp145;
	wire xformtmp136;
	assign xformtmp136 = in[57] | in[9];
	wire xformtmp129;
	assign xformtmp129 = xformtmp136 ^ in[65];
	wire xformtmp169;
	assign xformtmp169 = xformtmp139 | xformtmp129;
	wire xformtmp131;
	assign xformtmp131 = in[5] & xformtmp169;
	wire xformtmp171;
	assign xformtmp171 = xformtmp166 & xformtmp131;
	wire xformtmp138;
	assign xformtmp138 = in[131] ^ in[77];
	wire xformtmp137;
	assign xformtmp137 = xformtmp171 ^ xformtmp138;
	wire xformtmp134;
	assign xformtmp134 = xformtmp152 ^ xformtmp137;
	wire xformtmp167;
	assign xformtmp167 = in[99] ^ in[67];
	wire xformtmp159;
	assign xformtmp159 = in[0] & in[94];
	wire xformtmp128;
	assign xformtmp128 = xformtmp167 | xformtmp159;
	wire xformtmp161;
	assign xformtmp161 = xformtmp128 & in[48];
	wire xformtmp158;
	assign xformtmp158 = xformtmp161 & in[95];
	wire xformtmp160;
	assign xformtmp160 = in[73] | in[95];
	wire xformtmp165;
	assign xformtmp165 = in[38] | xformtmp160;
	wire xformtmp132;
	assign xformtmp132 = xformtmp158 & xformtmp165;
	wire xformtmp147;
	assign xformtmp147 = in[50] ^ in[8];
	wire xformtmp149;
	assign xformtmp149 = in[92] & in[98];
	wire xformtmp154;
	assign xformtmp154 = xformtmp147 & xformtmp149;
	wire xformtmp144;
	assign xformtmp144 = xformtmp132 & xformtmp154;
	assign out[3] = xformtmp134 | xformtmp144;
	assign out[4] = 1'b0;
	wire xformtmp175;
	assign xformtmp175 = in[118] & in[66];
	wire xformtmp177;
	assign xformtmp177 = in[66] | xformtmp175;
	wire xformtmp174;
	assign xformtmp174 = in[70] ^ xformtmp177;
	wire xformtmp176;
	assign xformtmp176 = in[66] & in[147];
	assign out[5] = xformtmp174 ^ xformtmp176;
	wire xformtmp178;
	assign xformtmp178 = in[22] | in[54];
	assign out[6] = xformtmp178 | in[84];
	assign out[78:7] = 72'b011010110110010101001100100100000101100001001000011001100011110011010100;
	assign out[79] = in[100];
endmodule

module tb();
    reg[79:0] results[1];
    reg[149:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%150b]", data[0]);
        #1
        $display("results = [%80b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
