module dut (out, in);
	output[29:0] out;
	input[49:0] in;
	wire origtmp1;
	wire origtmp2;
	wire origtmp3;
	wire origtmp4;
	wire origtmp5;
	wire origtmp6;
	wire origtmp7;
	wire origtmp8;
	wire origtmp9;
	wire origtmp10;
	wire origtmp11;
	wire origtmp12;
	wire origtmp13;
	wire origtmp14;
	wire origtmp15;
	wire origtmp16;
	wire origtmp17;
	wire origtmp18;
	wire origtmp19;
	wire origtmp20;
	wire origtmp21;
	wire origtmp22;
	wire origtmp23;
	wire origtmp24;
	wire origtmp25;
	wire origtmp26;
	wire origtmp27;
	wire origtmp28;
	wire origtmp29;
	wire origtmp30;
	wire origtmp31;
	wire origtmp32;
	wire origtmp33;
	wire origtmp34;
	wire origtmp35;
	wire origtmp36;
	wire origtmp37;
	wire origtmp38;
	wire origtmp39;
	wire origtmp40;
	wire origtmp41;
	wire origtmp42;
	wire origtmp43;
	wire origtmp44;
	wire origtmp45;
	wire origtmp46;
	wire origtmp47;
	wire origtmp48;
	wire origtmp49;
	wire origtmp50;
	wire origtmp51;
	wire origtmp52;
	wire origtmp53;
	wire origtmp54;
	wire origtmp55;
	wire origtmp56;
	wire origtmp57;
	wire origtmp58;
	wire origtmp59;
	wire origtmp60;
	wire origtmp61;
	wire origtmp62;
	wire origtmp63;
	wire origtmp64;
	wire origtmp65;
	wire origtmp66;
	wire origtmp67;
	wire origtmp68;
	wire origtmp69;
	wire origtmp70;
	wire origtmp71;
	wire origtmp72;
	assign out[10] = ~origtmp63;
	assign origtmp48 = origtmp31 | origtmp27;
	assign origtmp53 = in[41] & in[43];
	assign origtmp12 = origtmp51 | in[5];
	assign origtmp2 = in[32] ^ origtmp4;
	assign out[15] = origtmp65 ^ 1'b1;
	assign origtmp9 = in[42] | origtmp15;
	assign origtmp51 = origtmp49 & origtmp21;
	assign out[25] = ~1'b1;
	assign origtmp47 = in[28] & in[31];
	assign origtmp4 = ~origtmp6;
	assign out[7] = 1'b0 & 1'b1;
	assign origtmp41 = origtmp26 | origtmp22;
	assign origtmp34 = origtmp30 & in[16];
	assign origtmp32 = in[40];
	assign origtmp16 = in[24] | in[46];
	assign out[6] = ~origtmp62;
	assign origtmp17 = origtmp52 & origtmp10;
	assign origtmp18 = in[45] ^ origtmp37;
	assign origtmp5 = ~in[14];
	assign origtmp11 = origtmp29 & in[15];
	assign origtmp68 = ~1'b0;
	assign origtmp66 = 1'b0 ^ 1'b1;
	assign origtmp72 = in[2] ^ 1'b0;
	assign origtmp1 = origtmp2 | origtmp5;
	assign origtmp61 = in[3] | 1'b0;
	assign origtmp57 = origtmp59 | in[30];
	assign origtmp21 = origtmp39 & origtmp50;
	assign out[14] = ~1'b1;
	assign origtmp40 = in[39] | in[35];
	assign out[16] = 1'b0;
	assign origtmp45 = in[33] ^ in[47];
	assign origtmp15 = in[18] ^ origtmp23;
	assign origtmp54 = in[41] ^ in[21];
	assign origtmp62 = 1'b1 & 1'b0;
	assign origtmp39 = in[28] ^ origtmp35;
	assign origtmp69 = 1'b0 ^ 1'b0;
	assign origtmp67 = 1'b1;
	assign origtmp58 = in[36] ^ origtmp54;
	assign out[8] = 1'b1 & 1'b0;
	assign origtmp56 = origtmp57 | origtmp60;
	assign out[11] = 1'b1 ^ 1'b0;
	assign out[29] = 1'b1 ^ origtmp72;
	assign origtmp8 = origtmp11 & origtmp13;
	assign origtmp43 = origtmp24 & in[44];
	assign out[13] = ~1'b0;
	assign origtmp64 = 1'b0;
	assign origtmp49 = origtmp8 & origtmp44;
	assign out[4] = 1'b1 ^ 1'b0;
	assign origtmp25 = in[16] | origtmp9;
	assign origtmp10 = origtmp40 ^ origtmp38;
	assign out[2] = origtmp58 & origtmp56;
	assign origtmp52 = origtmp45 | in[49];
	assign origtmp7 = ~origtmp1;
	assign origtmp24 = origtmp19 | in[11];
	assign out[21] = origtmp68 & 1'b0;
	assign origtmp59 = in[26] ^ in[23];
	assign origtmp26 = origtmp33 & in[11];
	assign out[1] = origtmp17 & origtmp12;
	assign out[27] = origtmp70 ^ origtmp70;
	assign origtmp31 = origtmp25 | in[6];
	assign origtmp3 = in[20] | in[7];
	assign origtmp71 = 1'b1 ^ 1'b1;
	assign out[26] = 1'b1 ^ origtmp69;
	assign out[9] = 1'b1 | 1'b1;
	assign out[23] = 1'b1 ^ 1'b1;
	assign out[5] = ~1'b1;
	assign origtmp65 = 1'b0 | 1'b0;
	assign origtmp13 = origtmp14 | origtmp16;
	assign origtmp30 = origtmp48 | origtmp20;
	assign out[28] = origtmp71 | origtmp71;
	assign out[20] = origtmp67 | 1'b1;
	assign out[17] = origtmp66 & 1'b0;
	assign origtmp63 = 1'b1 ^ 1'b0;
	assign origtmp36 = in[17] | in[39];
	assign origtmp23 = in[22] ^ in[5];
	assign origtmp46 = in[1] ^ in[48];
	assign origtmp70 = ~1'b1;
	assign origtmp6 = in[14] ^ in[27];
	assign out[0] = origtmp7 ^ origtmp3;
	assign origtmp19 = in[34] ^ in[33];
	assign origtmp35 = in[0] | origtmp34;
	assign origtmp20 = ~origtmp47;
	assign origtmp42 = origtmp43 ^ in[37];
	assign origtmp55 = in[4] & in[8];
	assign origtmp44 = origtmp32 | origtmp46;
	assign origtmp60 = origtmp53 & origtmp55;
	assign origtmp33 = in[38] | origtmp36;
	assign out[3] = ~origtmp61;
	assign out[12] = 1'b1 | origtmp64;
	assign origtmp14 = in[22] & in[25];
	assign origtmp29 = in[19] & in[10];
	assign out[24] = 1'b1;
	assign origtmp27 = in[42] & in[12];
	assign out[18] = 1'b1 | 1'b1;
	assign out[22] = 1'b0 ^ 1'b1;
	assign origtmp50 = origtmp28 | origtmp42;
	assign out[19] = 1'b1 & 1'b0;
	assign origtmp38 = origtmp18 & in[13];
	assign origtmp37 = in[34] ^ in[35];
	assign origtmp28 = origtmp41 & in[48];
	assign origtmp22 = in[29] & in[9];
endmodule

module tb();
    reg[29:0] results[1];
    reg[49:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%50b]", data[0]);
        #1
        $display("results = [%30b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
