module dut (out, in);
	output[9:0] out;
	input[19:0] in;
	wire xformtemp30;
	wire xformtemp29;
	wire xformtemp28;
	wire xformtemp27;
	wire xformtemp26;
	wire xformtemp25;
	wire xformtemp24;
	wire xformtemp11;
	wire xformtemp10;
	wire xformtemp9;
	wire xformtemp8;
	wire xformtemp7;
	wire xformtemp6;
	wire xformtemp2;
	wire xformtemp1;
	wire xformtemp3;
	wire xformtemp4;
	wire xformtemp5;
	wire xformtemp12;
	wire xformtemp13;
	wire xformtemp14;
	wire xformtemp15;
	wire xformtemp16;
	wire xformtemp17;
	wire xformtemp18;
	wire xformtemp19;
	wire xformtemp20;
	wire xformtemp21;
	wire xformtemp22;
	wire xformtemp23;
	assign out[9] = xformtmp30 | in[8];
	assign out[8] = 1'b0;
	assign out[7] = 1'b0 & 1'b0;
	assign out[6] = 1'b0;
	assign out[5] = xformtmp29 & 1'b1;
	assign out[1] = xformtmp25 ^ in[1];
	assign out[0] = xformtmp3 ^ xformtmp19;
	assign out[2] = in[5] | xformtmp27;
	assign out[3] = in[19] | xformtmp28;
	assign out[4] = 1'b1;
	assign xformtmp30 = 1'b1;
	assign xformtmp29 = 1'b0 ^ 1'b0;
	assign xformtmp28 = in[19] ^ in[19];
	assign xformtmp27 = 1'b0;
	assign xformtmp26 = 1'b0 | in[1];
	assign xformtmp25 = xformtmp26 | xformtmp23;
	assign xformtmp24 = in[13] & in[12];
	assign xformtmp11 = xformtmp22 ^ xformtmp16;
	assign xformtmp10 = xformtmp20 | in[2];
	assign xformtmp9 = in[4] | xformtmp17;
	assign xformtmp8 = in[14] | in[3];
	assign xformtmp7 = in[11] & in[0];
	assign xformtmp6 = in[10] ^ in[15];
	assign xformtmp2 = in[17] | xformtmp10;
	assign xformtmp1 = xformtmp5 ^ in[6];
	assign xformtmp3 = xformtmp1 & xformtmp11;
	assign xformtmp4 = xformtmp14 ^ xformtmp15;
	assign xformtmp5 = in[2] | xformtmp9;
	assign xformtmp12 = xformtmp6 & in[6];
	assign xformtmp13 = in[17] & in[10];
	assign xformtmp14 = in[6] | in[16];
	assign xformtmp15 = xformtmp2 & xformtmp13;
	assign xformtmp16 = in[9] | xformtmp7;
	assign xformtmp17 = in[16] & 1'b1;
	assign xformtmp18 = xformtmp8 & 1'b1;
	assign xformtmp19 = xformtmp4 | xformtmp21;
	assign xformtmp20 = in[7] | in[10];
	assign xformtmp21 = xformtmp18 ^ in[4];
	assign xformtmp22 = xformtmp12 ^ in[7];
	assign xformtmp23 = in[18] | xformtmp24;
endmodule

module tb();
    reg[9:0] results[1];
    reg[19:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%20b]", data[0]);
        #1
        $display("results = [%10b]", results[0]);
        $writememb("results.txt", results);
    end 
endmodule
