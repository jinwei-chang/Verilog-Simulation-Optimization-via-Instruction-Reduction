module dut (out, in);
	output[499:0] out;
	input[1499:0] in;
	assign out[0] = in[544] | in[626];
	assign out[1] = 1'b1;
	assign out[2] = ~in[1456];
	assign out[3] = in[634] & in[1486];
	assign out[4] = in[735] & in[1344];
	assign out[6:5] = 2'b10;
	assign out[7] = in[383] & in[1474];
	assign out[11:8] = 4'b1011;
	assign out[12] = in[1366] | in[1379];
	assign out[14:13] = 2'b10;
	assign out[15] = in[749];
	assign out[18:16] = 3'b010;
	assign out[19] = in[905];
	assign out[20] = 1'b1;
	assign out[21] = in[817];
	assign out[22] = 1'b1;
	wire xformtmp59;
	assign xformtmp59 = in[330] | in[733];
	wire xformtmp60;
	assign xformtmp60 = ~xformtmp59;
	assign out[23] = in[330] ^ xformtmp60;
	assign out[24] = 1'b1;
	assign out[25] = ~in[952];
	assign out[29:26] = 4'b1000;
	assign out[30] = in[1139];
	assign out[31] = in[882];
	assign out[32] = in[123];
	assign out[38:33] = 6'b000010;
	assign out[39] = in[504];
	assign out[42:40] = 3'b000;
	assign out[43] = ~in[1416];
	assign out[44] = in[807] & in[1077];
	assign out[46:45] = 2'b10;
	assign out[47] = in[701] | in[870];
	assign out[48] = 1'b1;
	assign out[49] = in[83];
	assign out[52:50] = 3'b011;
	assign out[53] = in[106] & in[374];
	assign out[54] = ~in[953];
	assign out[56:55] = 2'b01;
	assign out[57] = ~in[1018];
	assign out[58] = in[1051];
	assign out[59] = in[289] | in[1336];
	assign out[60] = ~in[241];
	assign out[61] = ~in[812];
	assign out[62] = 1'b1;
	wire xformtmp2325;
	assign xformtmp2325 = ~in[516];
	assign out[63] = in[872] | xformtmp2325;
	assign out[64] = 1'b0;
	assign out[65] = in[320];
	assign out[68:66] = 3'b000;
	assign out[69] = ~in[166];
	assign out[80:70] = 11'b11100100010;
	assign out[81] = in[963];
	assign out[87:82] = 6'b010101;
	assign out[88] = in[1062] | in[1437];
	assign out[89] = 1'b0;
	assign out[90] = in[960] ^ in[1362];
	assign out[93:91] = 3'b100;
	wire xformtmp236;
	assign xformtmp236 = ~in[1074];
	assign out[94] = in[1357] | xformtmp236;
	assign out[95] = ~in[1293];
	assign out[97:96] = 2'b01;
	assign out[98] = in[585];
	assign out[100:99] = 2'b10;
	assign out[101] = in[1099] & in[1133];
	assign out[102] = 1'b0;
	wire xformtmp257;
	assign xformtmp257 = ~in[670];
	assign out[103] = in[1188] & xformtmp257;
	assign out[104] = in[851];
	assign out[107:105] = 3'b111;
	assign out[108] = in[387];
	assign out[111:109] = 3'b100;
	assign out[112] = in[461];
	assign out[114:113] = 2'b10;
	assign out[115] = in[1164];
	assign out[116] = in[1061] ^ in[1168];
	assign out[119:117] = 3'b010;
	assign out[120] = in[1417];
	assign out[121] = in[1402];
	assign out[124:122] = 3'b101;
	assign out[125] = in[98];
	assign out[126] = in[365];
	assign out[127] = ~in[1268];
	assign out[128] = 1'b1;
	assign out[129] = in[1241];
	assign out[135:130] = 6'b110100;
	assign out[136] = in[852] | in[1323];
	assign out[137] = in[1335];
	assign out[138] = 1'b0;
	assign out[139] = in[221] ^ in[1073];
	assign out[140] = in[228] & in[1044];
	assign out[141] = in[630];
	assign out[144:142] = 3'b011;
	wire xformtmp359;
	assign xformtmp359 = ~in[613];
	assign out[145] = in[420] ^ xformtmp359;
	assign out[146] = in[1143];
	assign out[148:147] = 2'b00;
	wire xformtmp367;
	assign xformtmp367 = in[828] ^ in[1387];
	wire xformtmp370;
	assign xformtmp370 = in[828] & in[1387];
	wire xformtmp371;
	assign xformtmp371 = ~xformtmp370;
	assign out[149] = xformtmp367 & xformtmp371;
	assign out[150] = in[1002];
	assign out[151] = 1'b0;
	assign out[152] = in[63] | in[847];
	assign out[153] = in[124] | in[1315];
	assign out[154] = in[384];
	assign out[155] = in[276];
	assign out[156] = ~in[9];
	assign out[157] = in[583] & in[709];
	assign out[158] = in[340] ^ in[545];
	assign out[159] = ~in[1167];
	assign out[164:160] = 5'b01111;
	assign out[165] = in[443] ^ in[1302];
	assign out[167:166] = 2'b11;
	assign out[168] = in[255] ^ in[510];
	assign out[169] = 1'b1;
	assign out[170] = ~in[35];
	assign out[171] = 1'b1;
	assign out[172] = in[82] & in[751];
	assign out[174:173] = 2'b01;
	assign out[175] = in[606];
	assign out[176] = 1'b1;
	wire xformtmp441;
	assign xformtmp441 = ~in[560];
	assign out[177] = in[97] & xformtmp441;
	assign out[180:178] = 3'b010;
	assign out[181] = in[115];
	assign out[183:182] = 2'b11;
	assign out[184] = in[185];
	assign out[185] = in[885];
	assign out[186] = in[715];
	assign out[187] = in[842];
	assign out[188] = in[501] | in[1269];
	assign out[189] = in[644];
	assign out[190] = 1'b1;
	assign out[191] = ~in[738];
	assign out[193:192] = 2'b10;
	assign out[194] = ~in[892];
	assign out[196:195] = 2'b11;
	assign out[197] = in[1243];
	assign out[198] = in[256];
	assign out[199] = 1'b1;
	assign out[200] = in[822];
	assign out[201] = in[222] & in[922];
	assign out[202] = in[1233];
	assign out[203] = ~in[800];
	assign out[204] = in[480] ^ in[1240];
	assign out[205] = 1'b0;
	assign out[206] = in[1394];
	assign out[207] = 1'b1;
	assign out[208] = in[894] | in[1255];
	assign out[209] = 1'b1;
	assign out[210] = in[137] ^ in[1152];
	assign out[212:211] = 2'b01;
	wire xformtmp525;
	assign xformtmp525 = in[422] | in[891];
	assign out[213] = ~xformtmp525;
	wire xformtmp528;
	assign xformtmp528 = ~in[1414];
	wire xformtmp530;
	assign xformtmp530 = in[920] ^ in[1414];
	assign out[214] = xformtmp528 | xformtmp530;
	wire xformtmp531;
	assign xformtmp531 = ~in[339];
	wire xformtmp532;
	assign xformtmp532 = in[203] & xformtmp531;
	assign out[215] = ~xformtmp532;
	assign out[219:216] = 4'b1110;
	assign out[220] = in[488] & in[721];
	assign out[221] = in[479];
	assign out[224:222] = 3'b000;
	assign out[225] = ~in[99];
	assign out[226] = 1'b0;
	assign out[227] = in[411] & in[1060];
	assign out[230:228] = 3'b001;
	assign out[231] = ~in[152];
	assign out[232] = 1'b1;
	assign out[233] = in[451] & in[519];
	assign out[234] = in[10] | in[201];
	assign out[235] = 1'b0;
	assign out[236] = in[1272];
	assign out[240:237] = 4'b1100;
	assign out[241] = ~in[1393];
	assign out[251:242] = 10'b1100000011;
	wire xformtmp628;
	assign xformtmp628 = ~in[838];
	wire xformtmp629;
	assign xformtmp629 = ~in[1460];
	assign out[252] = xformtmp628 | xformtmp629;
	assign out[253] = in[380] | in[1479];
	assign out[254] = 1'b0;
	assign out[255] = in[503];
	wire xformtmp635;
	assign xformtmp635 = ~in[368];
	wire xformtmp634;
	assign xformtmp634 = in[130] & xformtmp635;
	wire xformtmp636;
	assign xformtmp636 = ~in[130];
	assign out[256] = xformtmp634 ^ xformtmp636;
	assign out[257] = 1'b1;
	wire xformtmp640;
	assign xformtmp640 = ~in[364];
	assign out[258] = in[7] | xformtmp640;
	assign out[259] = in[1345] | in[1495];
	assign out[261:260] = 2'b10;
	assign out[262] = ~in[593];
	assign out[264:263] = 2'b01;
	assign out[265] = in[431];
	assign out[268:266] = 3'b011;
	assign out[269] = in[162] | in[1100];
	assign out[271:270] = 2'b10;
	assign out[272] = ~in[207];
	assign out[275:273] = 3'b010;
	assign out[276] = in[275] & in[1021];
	wire xformtmp2311;
	assign xformtmp2311 = ~in[1157];
	assign out[277] = in[976] & xformtmp2311;
	assign out[278] = in[757];
	assign out[279] = in[862];
	assign out[280] = 1'b1;
	assign out[281] = in[977] | in[1257];
	assign out[284:282] = 3'b001;
	assign out[285] = ~in[534];
	wire xformtmp724;
	assign xformtmp724 = ~in[208];
	wire xformtmp725;
	assign xformtmp725 = in[220] ^ xformtmp724;
	assign out[286] = ~xformtmp725;
	wire xformtmp728;
	assign xformtmp728 = ~in[388];
	assign out[287] = in[274] | xformtmp728;
	assign out[288] = 1'b1;
	assign out[289] = in[767];
	assign out[290] = ~in[1227];
	assign out[291] = ~in[500];
	assign out[293:292] = 2'b11;
	assign out[294] = in[235] ^ in[944];
	assign out[295] = 1'b1;
	assign out[296] = in[1329];
	assign out[297] = 1'b0;
	assign out[298] = in[614];
	assign out[300:299] = 2'b10;
	assign out[301] = in[1171];
	assign out[303:302] = 2'b00;
	assign out[304] = ~in[695];
	assign out[305] = ~in[784];
	assign out[306] = ~in[884];
	assign out[307] = in[1230] | in[1435];
	assign out[308] = 1'b0;
	assign out[309] = in[257] ^ in[399];
	wire xformtmp2371;
	assign xformtmp2371 = in[810] & in[1179];
	assign out[310] = ~xformtmp2371;
	assign out[311] = 1'b1;
	assign out[312] = in[108] ^ in[502];
	assign out[314:313] = 2'b00;
	assign out[315] = in[55] & in[1489];
	assign out[323:316] = 8'b00010110;
	wire xformtmp806;
	assign xformtmp806 = ~in[464];
	assign out[324] = in[492] & xformtmp806;
	assign out[326:325] = 2'b01;
	wire xformtmp812;
	assign xformtmp812 = ~in[991];
	assign out[327] = in[1332] ^ xformtmp812;
	assign out[329:328] = 2'b10;
	assign out[330] = in[341] | in[432];
	assign out[331] = ~in[1458];
	assign out[337:332] = 6'b001110;
	assign out[338] = in[640];
	assign out[342:339] = 4'b1001;
	assign out[343] = in[651] ^ in[825];
	assign out[344] = ~in[491];
	assign out[345] = ~in[425];
	assign out[346] = in[138];
	assign out[347] = in[298] & in[926];
	assign out[348] = in[148];
	assign out[349] = in[70];
	assign out[351:350] = 2'b00;
	assign out[352] = in[486] & in[1395];
	assign out[353] = 1'b0;
	assign out[354] = in[286] | in[297];
	assign out[355] = 1'b1;
	assign out[356] = in[2] & in[96];
	assign out[358:357] = 2'b10;
	wire xformtmp894;
	assign xformtmp894 = in[804] ^ in[1447];
	wire xformtmp895;
	assign xformtmp895 = in[804] | in[1447];
	assign out[359] = xformtmp894 & xformtmp895;
	assign out[362:360] = 3'b001;
	assign out[363] = in[270] & in[468];
	assign out[364] = 1'b1;
	assign out[365] = in[829] ^ in[1138];
	wire xformtmp905;
	assign xformtmp905 = ~in[29];
	assign out[366] = in[1134] & xformtmp905;
	assign out[367] = 1'b0;
	assign out[368] = in[386] & in[589];
	assign out[369] = ~in[316];
	assign out[374:370] = 5'b00111;
	assign out[375] = in[116] ^ in[780];
	assign out[376] = in[478];
	assign out[378:377] = 2'b00;
	assign out[379] = in[436];
	assign out[381:380] = 2'b10;
	assign out[382] = ~in[347];
	assign out[383] = in[1350];
	assign out[384] = in[318] & in[931];
	assign out[388:385] = 4'b0111;
	assign out[389] = in[1271];
	assign out[390] = in[105] & in[874];
	assign out[391] = 1'b1;
	wire xformtmp969;
	assign xformtmp969 = ~in[704];
	assign out[392] = in[567] & xformtmp969;
	assign out[393] = in[536];
	assign out[394] = 1'b1;
	assign out[395] = in[446] ^ in[1039];
	assign out[397:396] = 2'b00;
	assign out[398] = in[1413];
	assign out[399] = in[412];
	assign out[400] = in[1020];
	wire xformtmp994;
	assign xformtmp994 = ~in[53];
	assign out[401] = in[1106] & xformtmp994;
	wire xformtmp996;
	assign xformtmp996 = ~in[47];
	assign out[402] = in[1169] & xformtmp996;
	assign out[403] = in[1064];
	assign out[404] = 1'b0;
	assign out[405] = in[602];
	assign out[409:406] = 4'b1101;
	assign out[410] = in[77] & in[1462];
	assign out[411] = in[802];
	assign out[412] = 1'b0;
	assign out[413] = in[72];
	assign out[416:414] = 3'b100;
	assign out[417] = in[1289];
	assign out[418] = 1'b1;
	assign out[419] = in[1123];
	assign out[420] = 1'b1;
	assign out[421] = in[1311];
	assign out[422] = 1'b0;
	assign out[423] = in[816];
	assign out[426:424] = 3'b001;
	assign out[427] = in[369] & in[1423];
	assign out[428] = in[726] ^ in[938];
	assign out[434:429] = 6'b101100;
	assign out[435] = in[896];
	assign out[438:436] = 3'b000;
	assign out[439] = in[1178];
	assign out[441:440] = 2'b00;
	wire xformtmp1097;
	assign xformtmp1097 = ~in[582];
	assign out[442] = in[898] | xformtmp1097;
	assign out[443] = in[1258];
	assign out[444] = ~in[1047];
	assign out[448:445] = 4'b0101;
	assign out[449] = in[541];
	assign out[450] = in[273];
	assign out[452:451] = 2'b10;
	wire xformtmp1132;
	assign xformtmp1132 = ~in[818];
	assign out[453] = in[90] & xformtmp1132;
	assign out[454] = ~in[1383];
	assign out[455] = ~in[188];
	assign out[456] = in[328];
	assign out[457] = 1'b0;
	assign out[458] = in[653];
	assign out[460:459] = 2'b00;
	assign out[461] = in[252];
	assign out[462] = 1'b0;
	assign out[463] = in[554];
	assign out[464] = 1'b0;
	assign out[465] = in[787];
	assign out[466] = in[366];
	assign out[467] = ~in[1246];
	assign out[468] = 1'b1;
	assign out[469] = in[600];
	assign out[474:470] = 5'b10110;
	assign out[475] = in[332];
	assign out[476] = in[557] ^ in[1239];
	assign out[477] = ~in[110];
	assign out[479:478] = 2'b10;
	assign out[480] = in[1298] & in[1497];
	assign out[482:481] = 2'b10;
	wire xformtmp2339;
	assign xformtmp2339 = in[649] ^ in[1400];
	wire xformtmp1211;
	assign xformtmp1211 = in[649] | in[1400];
	wire xformtmp1213;
	assign xformtmp1213 = xformtmp2339 | xformtmp1211;
	assign out[483] = xformtmp1213 ^ xformtmp2339;
	assign out[484] = ~in[564];
	assign out[485] = in[338] ^ in[1339];
	assign out[486] = in[927] & in[1204];
	assign out[490:487] = 4'b0001;
	assign out[491] = in[294] ^ in[1141];
	assign out[492] = ~in[79];
	assign out[493] = 1'b0;
	assign out[494] = in[627];
	assign out[495] = 1'b1;
	assign out[496] = in[136];
	assign out[497] = 1'b0;
	wire xformtmp2275;
	assign xformtmp2275 = ~in[474];
	assign out[498] = in[972] & xformtmp2275;
	wire xformtmp1602;
	assign xformtmp1602 = in[518] | in[1042];
	wire xformtmp2076;
	assign xformtmp2076 = in[830] | xformtmp1602;
	wire xformtmp1636;
	assign xformtmp1636 = in[52] | in[785];
	wire xformtmp1356;
	assign xformtmp1356 = in[457] ^ in[1494];
	wire xformtmp1421;
	assign xformtmp1421 = in[605] ^ xformtmp1356;
	wire xformtmp2027;
	assign xformtmp2027 = in[584] ^ in[883];
	wire xformtmp1892;
	assign xformtmp1892 = xformtmp1421 & xformtmp2027;
	wire xformtmp1771;
	assign xformtmp1771 = in[694] & xformtmp1892;
	wire xformtmp1925;
	assign xformtmp1925 = in[890] ^ xformtmp1771;
	wire xformtmp1375;
	assign xformtmp1375 = xformtmp1636 ^ xformtmp1925;
	wire xformtmp1811;
	assign xformtmp1811 = in[158] ^ in[327];
	wire xformtmp1542;
	assign xformtmp1542 = in[392] | xformtmp1811;
	wire xformtmp1785;
	assign xformtmp1785 = in[489] | in[759];
	wire xformtmp2109;
	assign xformtmp2109 = xformtmp1542 ^ xformtmp1785;
	wire xformtmp1336;
	assign xformtmp1336 = in[1028] | xformtmp2109;
	wire xformtmp1397;
	assign xformtmp1397 = in[21] ^ in[811];
	wire xformtmp2043;
	assign xformtmp2043 = in[1409] ^ xformtmp1397;
	wire xformtmp1337;
	assign xformtmp1337 = in[1029] | xformtmp2043;
	wire xformtmp2079;
	assign xformtmp2079 = xformtmp1336 ^ xformtmp1337;
	wire xformtmp1635;
	assign xformtmp1635 = in[542] | xformtmp2079;
	wire xformtmp1997;
	assign xformtmp1997 = in[1220] ^ in[1373];
	wire xformtmp1298;
	assign xformtmp1298 = in[543] | xformtmp1997;
	wire xformtmp1475;
	assign xformtmp1475 = in[897] ^ in[1212];
	wire xformtmp1596;
	assign xformtmp1596 = in[209] | in[1122];
	wire xformtmp1610;
	assign xformtmp1610 = xformtmp1475 & xformtmp1596;
	wire xformtmp2211;
	assign xformtmp2211 = in[1312] | xformtmp1610;
	wire xformtmp1871;
	assign xformtmp1871 = in[413] | in[591];
	wire xformtmp2229;
	assign xformtmp2229 = in[1292] | xformtmp1871;
	wire xformtmp1934;
	assign xformtmp1934 = xformtmp2211 & xformtmp2229;
	wire xformtmp1783;
	assign xformtmp1783 = xformtmp1298 ^ xformtmp1934;
	wire xformtmp1710;
	assign xformtmp1710 = in[601] & xformtmp1783;
	wire xformtmp1676;
	assign xformtmp1676 = xformtmp1635 | xformtmp1710;
	wire xformtmp1913;
	assign xformtmp1913 = xformtmp1375 ^ xformtmp1676;
	wire xformtmp1851;
	assign xformtmp1851 = in[36] & in[669];
	wire xformtmp1889;
	assign xformtmp1889 = in[752] ^ in[758];
	wire xformtmp1248;
	assign xformtmp1248 = in[1173] ^ xformtmp1889;
	wire xformtmp1998;
	assign xformtmp1998 = in[303] & in[1248];
	wire xformtmp2103;
	assign xformtmp2103 = in[921] & xformtmp1998;
	wire xformtmp1410;
	assign xformtmp1410 = xformtmp1248 ^ xformtmp2103;
	wire xformtmp1246;
	assign xformtmp1246 = in[903] | xformtmp1410;
	wire xformtmp1510;
	assign xformtmp1510 = in[193] ^ in[301];
	wire xformtmp1315;
	assign xformtmp1315 = in[119] | in[1033];
	wire xformtmp1545;
	assign xformtmp1545 = in[1190] ^ in[1310];
	wire xformtmp1825;
	assign xformtmp1825 = in[992] ^ xformtmp1545;
	wire xformtmp2141;
	assign xformtmp2141 = in[248] | in[1434];
	wire xformtmp1970;
	assign xformtmp1970 = xformtmp1825 ^ xformtmp2141;
	wire xformtmp2254;
	assign xformtmp2254 = xformtmp1315 & xformtmp1970;
	wire xformtmp2150;
	assign xformtmp2150 = xformtmp1510 | xformtmp2254;
	wire xformtmp2224;
	assign xformtmp2224 = xformtmp1246 ^ xformtmp2150;
	wire xformtmp1299;
	assign xformtmp1299 = xformtmp1851 ^ xformtmp2224;
	wire xformtmp1436;
	assign xformtmp1436 = in[750] | in[1286];
	wire xformtmp1843;
	assign xformtmp1843 = in[172] | xformtmp1436;
	wire xformtmp1942;
	assign xformtmp1942 = in[1451] | xformtmp1843;
	wire xformtmp1668;
	assign xformtmp1668 = in[512] | xformtmp1942;
	wire xformtmp2232;
	assign xformtmp2232 = in[473] & in[714];
	wire xformtmp1517;
	assign xformtmp1517 = in[1305] ^ xformtmp2232;
	wire xformtmp2125;
	assign xformtmp2125 = in[561] | xformtmp1517;
	wire xformtmp2095;
	assign xformtmp2095 = in[1147] | xformtmp2125;
	wire xformtmp1694;
	assign xformtmp1694 = xformtmp1668 & xformtmp2095;
	wire xformtmp1908;
	assign xformtmp1908 = in[64] ^ in[1322];
	wire xformtmp1685;
	assign xformtmp1685 = in[575] ^ xformtmp1908;
	wire xformtmp1626;
	assign xformtmp1626 = in[1472] ^ xformtmp1685;
	wire xformtmp1977;
	assign xformtmp1977 = in[406] & xformtmp1626;
	wire xformtmp2046;
	assign xformtmp2046 = in[959] & xformtmp1977;
	wire xformtmp1525;
	assign xformtmp1525 = xformtmp1694 | xformtmp2046;
	wire xformtmp1706;
	assign xformtmp1706 = xformtmp1299 | xformtmp1525;
	wire xformtmp1651;
	assign xformtmp1651 = in[756] & in[1213];
	wire xformtmp1283;
	assign xformtmp1283 = in[1022] ^ xformtmp1651;
	wire xformtmp2165;
	assign xformtmp2165 = in[81] ^ xformtmp1283;
	wire xformtmp1573;
	assign xformtmp1573 = xformtmp1706 | xformtmp2165;
	wire xformtmp1322;
	assign xformtmp1322 = in[344] ^ in[535];
	wire xformtmp1473;
	assign xformtmp1473 = in[762] & in[1026];
	wire xformtmp1632;
	assign xformtmp1632 = xformtmp1322 ^ xformtmp1473;
	wire xformtmp1404;
	assign xformtmp1404 = in[1237] & in[1277];
	wire xformtmp1455;
	assign xformtmp1455 = in[1438] & xformtmp1404;
	wire xformtmp1659;
	assign xformtmp1659 = in[34] | in[281];
	wire xformtmp2190;
	assign xformtmp2190 = xformtmp1455 | xformtmp1659;
	wire xformtmp1841;
	assign xformtmp1841 = in[1014] & xformtmp2190;
	wire xformtmp1569;
	assign xformtmp1569 = xformtmp1632 ^ xformtmp1841;
	wire xformtmp1605;
	assign xformtmp1605 = in[659] | in[771];
	wire xformtmp1485;
	assign xformtmp1485 = in[28] & in[452];
	wire xformtmp2024;
	assign xformtmp2024 = in[1367] ^ xformtmp1485;
	wire xformtmp1682;
	assign xformtmp1682 = in[129] | xformtmp2024;
	wire xformtmp2000;
	assign xformtmp2000 = in[293] ^ xformtmp1682;
	wire xformtmp2202;
	assign xformtmp2202 = in[126] ^ xformtmp2000;
	wire xformtmp2006;
	assign xformtmp2006 = xformtmp1605 ^ xformtmp2202;
	wire xformtmp2161;
	assign xformtmp2161 = in[1158] | in[1436];
	wire xformtmp2158;
	assign xformtmp2158 = in[15] ^ xformtmp2161;
	wire xformtmp1989;
	assign xformtmp1989 = xformtmp2006 ^ xformtmp2158;
	wire xformtmp1929;
	assign xformtmp1929 = in[857] & xformtmp1989;
	wire xformtmp2157;
	assign xformtmp2157 = xformtmp1569 | xformtmp1929;
	wire xformtmp1677;
	assign xformtmp1677 = xformtmp1573 | xformtmp2157;
	wire xformtmp1311;
	assign xformtmp1311 = in[571] ^ in[1072];
	wire xformtmp1371;
	assign xformtmp1371 = in[1121] | xformtmp1311;
	wire xformtmp1429;
	assign xformtmp1429 = in[211] & in[378];
	wire xformtmp1449;
	assign xformtmp1449 = in[1] & in[1485];
	wire xformtmp1725;
	assign xformtmp1725 = in[23] & in[525];
	wire xformtmp1291;
	assign xformtmp1291 = xformtmp1449 & xformtmp1725;
	wire xformtmp1844;
	assign xformtmp1844 = in[652] & in[982];
	wire xformtmp1259;
	assign xformtmp1259 = in[441] ^ in[533];
	wire xformtmp2177;
	assign xformtmp2177 = in[213] ^ xformtmp1259;
	wire xformtmp2212;
	assign xformtmp2212 = xformtmp1844 ^ xformtmp2177;
	wire xformtmp1509;
	assign xformtmp1509 = xformtmp1291 & xformtmp2212;
	wire xformtmp1695;
	assign xformtmp1695 = xformtmp1429 | xformtmp1509;
	wire xformtmp1546;
	assign xformtmp1546 = xformtmp1371 & xformtmp1695;
	wire xformtmp1806;
	assign xformtmp1806 = in[624] ^ in[1333];
	wire xformtmp1810;
	assign xformtmp1810 = in[282] | xformtmp1806;
	wire xformtmp1631;
	assign xformtmp1631 = in[620] & in[1174];
	wire xformtmp1269;
	assign xformtmp1269 = in[1109] | xformtmp1631;
	wire xformtmp1689;
	assign xformtmp1689 = in[766] ^ in[948];
	wire xformtmp1697;
	assign xformtmp1697 = in[508] & xformtmp1689;
	wire xformtmp2110;
	assign xformtmp2110 = xformtmp1269 | xformtmp1697;
	wire xformtmp1923;
	assign xformtmp1923 = xformtmp1810 & xformtmp2110;
	wire xformtmp1331;
	assign xformtmp1331 = in[763] | in[1369];
	wire xformtmp2057;
	assign xformtmp2057 = in[955] ^ xformtmp1331;
	wire xformtmp1261;
	assign xformtmp1261 = xformtmp1923 & xformtmp2057;
	wire xformtmp1661;
	assign xformtmp1661 = in[1353] | in[1404];
	wire xformtmp1590;
	assign xformtmp1590 = in[358] ^ in[1313];
	wire xformtmp1708;
	assign xformtmp1708 = in[866] | in[1471];
	wire xformtmp1633;
	assign xformtmp1633 = in[456] & xformtmp1708;
	wire xformtmp2048;
	assign xformtmp2048 = in[149] | in[173];
	wire xformtmp1561;
	assign xformtmp1561 = xformtmp1633 | xformtmp2048;
	wire xformtmp1876;
	assign xformtmp1876 = in[1275] & xformtmp1561;
	wire xformtmp1669;
	assign xformtmp1669 = xformtmp1590 & xformtmp1876;
	wire xformtmp1355;
	assign xformtmp1355 = xformtmp1661 | xformtmp1669;
	wire xformtmp1251;
	assign xformtmp1251 = xformtmp1261 | xformtmp1355;
	wire xformtmp1621;
	assign xformtmp1621 = in[135] ^ in[176];
	wire xformtmp1407;
	assign xformtmp1407 = in[966] & xformtmp1621;
	wire xformtmp1705;
	assign xformtmp1705 = xformtmp1251 ^ xformtmp1407;
	wire xformtmp1411;
	assign xformtmp1411 = xformtmp1546 | xformtmp1705;
	wire xformtmp1946;
	assign xformtmp1946 = in[604] & in[720];
	wire xformtmp1738;
	assign xformtmp1738 = in[1465] | xformtmp1946;
	wire xformtmp2155;
	assign xformtmp2155 = in[5] | in[1201];
	wire xformtmp1630;
	assign xformtmp1630 = xformtmp1738 | xformtmp2155;
	wire xformtmp1797;
	assign xformtmp1797 = in[322] & in[1048];
	wire xformtmp1665;
	assign xformtmp1665 = in[980] ^ xformtmp1797;
	wire xformtmp1937;
	assign xformtmp1937 = in[498] ^ xformtmp1665;
	wire xformtmp1647;
	assign xformtmp1647 = in[529] | xformtmp1937;
	wire xformtmp1678;
	assign xformtmp1678 = xformtmp1630 & xformtmp1647;
	wire xformtmp1687;
	assign xformtmp1687 = in[1408] | in[1475];
	wire xformtmp1719;
	assign xformtmp1719 = in[1380] ^ xformtmp1687;
	wire xformtmp2070;
	assign xformtmp2070 = in[62] & in[731];
	wire xformtmp2086;
	assign xformtmp2086 = xformtmp1719 & xformtmp2070;
	wire xformtmp2204;
	assign xformtmp2204 = xformtmp1678 & xformtmp2086;
	wire xformtmp1723;
	assign xformtmp1723 = xformtmp1411 | xformtmp2204;
	wire xformtmp2061;
	assign xformtmp2061 = xformtmp1677 | xformtmp1723;
	wire xformtmp2192;
	assign xformtmp2192 = xformtmp1913 & xformtmp2061;
	wire xformtmp1279;
	assign xformtmp1279 = xformtmp2076 | xformtmp2192;
	wire xformtmp1779;
	assign xformtmp1779 = in[227] ^ in[1419];
	wire xformtmp1987;
	assign xformtmp1987 = in[770] | xformtmp1779;
	wire xformtmp1657;
	assign xformtmp1657 = in[530] | xformtmp1987;
	wire xformtmp1566;
	assign xformtmp1566 = in[1244] & in[1378];
	wire xformtmp1753;
	assign xformtmp1753 = in[237] | in[913];
	wire xformtmp1615;
	assign xformtmp1615 = in[599] ^ xformtmp1753;
	wire xformtmp1571;
	assign xformtmp1571 = in[983] & xformtmp1615;
	wire xformtmp1419;
	assign xformtmp1419 = xformtmp1566 ^ xformtmp1571;
	wire xformtmp1412;
	assign xformtmp1412 = in[381] ^ in[581];
	wire xformtmp1389;
	assign xformtmp1389 = in[742] | xformtmp1412;
	wire xformtmp1653;
	assign xformtmp1653 = in[837] ^ xformtmp1389;
	wire xformtmp2092;
	assign xformtmp2092 = xformtmp1419 | xformtmp1653;
	wire xformtmp1567;
	assign xformtmp1567 = in[472] | xformtmp2092;
	wire xformtmp1272;
	assign xformtmp1272 = in[41] | xformtmp1567;
	wire xformtmp1805;
	assign xformtmp1805 = in[164] | in[1036];
	wire xformtmp1820;
	assign xformtmp1820 = in[427] ^ xformtmp1805;
	wire xformtmp1264;
	assign xformtmp1264 = in[1294] ^ xformtmp1820;
	wire xformtmp1862;
	assign xformtmp1862 = in[300] & in[314];
	wire xformtmp1384;
	assign xformtmp1384 = in[879] | xformtmp1862;
	wire xformtmp1376;
	assign xformtmp1376 = in[462] ^ xformtmp1384;
	wire xformtmp1921;
	assign xformtmp1921 = in[645] & in[813];
	wire xformtmp1927;
	assign xformtmp1927 = in[251] & in[460];
	wire xformtmp1833;
	assign xformtmp1833 = xformtmp1921 & xformtmp1927;
	wire xformtmp1570;
	assign xformtmp1570 = xformtmp1376 | xformtmp1833;
	wire xformtmp2044;
	assign xformtmp2044 = xformtmp1264 & xformtmp1570;
	wire xformtmp1848;
	assign xformtmp1848 = xformtmp1272 ^ xformtmp2044;
	wire xformtmp1991;
	assign xformtmp1991 = xformtmp1657 & xformtmp1848;
	wire xformtmp1365;
	assign xformtmp1365 = xformtmp1279 & xformtmp1991;
	wire xformtmp1274;
	assign xformtmp1274 = in[377] | in[612];
	wire xformtmp1402;
	assign xformtmp1402 = in[970] | in[1013];
	wire xformtmp2036;
	assign xformtmp2036 = in[93] | xformtmp1402;
	wire xformtmp1838;
	assign xformtmp1838 = xformtmp1274 & xformtmp2036;
	wire xformtmp1538;
	assign xformtmp1538 = xformtmp1365 | xformtmp1838;
	wire xformtmp1645;
	assign xformtmp1645 = in[820] ^ in[1499];
	wire xformtmp2054;
	assign xformtmp2054 = in[89] & xformtmp1645;
	wire xformtmp1704;
	assign xformtmp1704 = in[867] & xformtmp2054;
	wire xformtmp1413;
	assign xformtmp1413 = in[56] & in[1217];
	wire xformtmp2028;
	assign xformtmp2028 = in[531] | xformtmp1413;
	wire xformtmp2089;
	assign xformtmp2089 = in[362] & in[375];
	wire xformtmp1378;
	assign xformtmp1378 = xformtmp2028 | xformtmp2089;
	wire xformtmp1886;
	assign xformtmp1886 = in[710] | in[899];
	wire xformtmp1735;
	assign xformtmp1735 = in[917] | xformtmp1886;
	wire xformtmp1814;
	assign xformtmp1814 = in[943] | xformtmp1735;
	wire xformtmp2115;
	assign xformtmp2115 = in[1348] ^ xformtmp1814;
	wire xformtmp2180;
	assign xformtmp2180 = in[1124] ^ xformtmp2115;
	wire xformtmp1887;
	assign xformtmp1887 = xformtmp1378 | xformtmp2180;
	wire xformtmp2059;
	assign xformtmp2059 = in[777] | in[1131];
	wire xformtmp1574;
	assign xformtmp1574 = in[396] | xformtmp2059;
	wire xformtmp2153;
	assign xformtmp2153 = in[1291] | xformtmp1574;
	wire xformtmp2210;
	assign xformtmp2210 = in[1488] | xformtmp2153;
	wire xformtmp2010;
	assign xformtmp2010 = xformtmp1887 ^ xformtmp2210;
	wire xformtmp2183;
	assign xformtmp2183 = in[621] & in[1087];
	wire xformtmp1736;
	assign xformtmp1736 = in[779] | xformtmp2183;
	wire xformtmp1463;
	assign xformtmp1463 = in[402] ^ xformtmp1736;
	wire xformtmp2167;
	assign xformtmp2167 = in[428] ^ in[1228];
	wire xformtmp1576;
	assign xformtmp1576 = in[836] | xformtmp2167;
	wire xformtmp1739;
	assign xformtmp1739 = xformtmp1463 | xformtmp1576;
	wire xformtmp2025;
	assign xformtmp2025 = in[741] | xformtmp1739;
	wire xformtmp1250;
	assign xformtmp1250 = in[691] | in[1477];
	wire xformtmp1484;
	assign xformtmp1484 = in[400] & in[1478];
	wire xformtmp1718;
	assign xformtmp1718 = in[1024] | xformtmp1484;
	wire xformtmp1874;
	assign xformtmp1874 = xformtmp1250 | xformtmp1718;
	wire xformtmp2236;
	assign xformtmp2236 = in[665] & xformtmp1874;
	wire xformtmp2071;
	assign xformtmp2071 = xformtmp2025 ^ xformtmp2236;
	wire xformtmp2213;
	assign xformtmp2213 = xformtmp2010 & xformtmp2071;
	wire xformtmp1768;
	assign xformtmp1768 = xformtmp1704 | xformtmp2213;
	wire xformtmp2069;
	assign xformtmp2069 = in[1082] ^ in[1491];
	wire xformtmp1335;
	assign xformtmp1335 = in[1266] & xformtmp2069;
	wire xformtmp1903;
	assign xformtmp1903 = in[734] ^ in[941];
	wire xformtmp1673;
	assign xformtmp1673 = in[985] | xformtmp1903;
	wire xformtmp1346;
	assign xformtmp1346 = xformtmp1335 ^ xformtmp1673;
	wire xformtmp1535;
	assign xformtmp1535 = in[0] ^ in[409];
	wire xformtmp1363;
	assign xformtmp1363 = in[66] | xformtmp1535;
	wire xformtmp1293;
	assign xformtmp1293 = in[225] | xformtmp1363;
	wire xformtmp1252;
	assign xformtmp1252 = in[654] ^ in[964];
	wire xformtmp2175;
	assign xformtmp2175 = in[1035] ^ xformtmp1252;
	wire xformtmp1625;
	assign xformtmp1625 = xformtmp1293 & xformtmp2175;
	wire xformtmp1275;
	assign xformtmp1275 = in[1095] ^ in[1464];
	wire xformtmp1324;
	assign xformtmp1324 = in[1187] & xformtmp1275;
	wire xformtmp1592;
	assign xformtmp1592 = in[1215] ^ xformtmp1324;
	wire xformtmp1740;
	assign xformtmp1740 = in[598] | in[1037];
	wire xformtmp1786;
	assign xformtmp1786 = in[38] & xformtmp1740;
	wire xformtmp1310;
	assign xformtmp1310 = in[429] ^ in[860];
	wire xformtmp1467;
	assign xformtmp1467 = in[625] & in[679];
	wire xformtmp2085;
	assign xformtmp2085 = xformtmp1310 | xformtmp1467;
	wire xformtmp1373;
	assign xformtmp1373 = in[1205] ^ xformtmp2085;
	wire xformtmp2077;
	assign xformtmp2077 = in[447] & in[1411];
	wire xformtmp1932;
	assign xformtmp1932 = in[662] & in[1025];
	wire xformtmp2090;
	assign xformtmp2090 = in[910] ^ xformtmp1932;
	wire xformtmp1722;
	assign xformtmp1722 = xformtmp2077 | xformtmp2090;
	wire xformtmp1472;
	assign xformtmp1472 = xformtmp1373 | xformtmp1722;
	wire xformtmp1856;
	assign xformtmp1856 = in[199] | in[725];
	wire xformtmp1350;
	assign xformtmp1350 = in[397] ^ xformtmp1856;
	wire xformtmp1796;
	assign xformtmp1796 = in[1016] & in[1110];
	wire xformtmp2174;
	assign xformtmp2174 = xformtmp1350 ^ xformtmp1796;
	wire xformtmp1593;
	assign xformtmp1593 = in[635] | xformtmp2174;
	wire xformtmp2100;
	assign xformtmp2100 = xformtmp1472 | xformtmp1593;
	wire xformtmp1641;
	assign xformtmp1641 = xformtmp1786 & xformtmp2100;
	wire xformtmp1791;
	assign xformtmp1791 = xformtmp1592 & xformtmp1641;
	wire xformtmp1415;
	assign xformtmp1415 = xformtmp1625 | xformtmp1791;
	wire xformtmp2118;
	assign xformtmp2118 = xformtmp1346 | xformtmp1415;
	wire xformtmp1441;
	assign xformtmp1441 = xformtmp1768 | xformtmp2118;
	wire xformtmp1734;
	assign xformtmp1734 = in[1065] ^ in[1466];
	wire xformtmp1660;
	assign xformtmp1660 = in[1091] ^ xformtmp1734;
	wire xformtmp1563;
	assign xformtmp1563 = in[348] | in[703];
	wire xformtmp1650;
	assign xformtmp1650 = in[935] ^ xformtmp1563;
	wire xformtmp1952;
	assign xformtmp1952 = in[597] & in[1092];
	wire xformtmp1386;
	assign xformtmp1386 = xformtmp1650 & xformtmp1952;
	wire xformtmp1242;
	assign xformtmp1242 = in[65] ^ in[1385];
	wire xformtmp1495;
	assign xformtmp1495 = in[1090] | xformtmp1242;
	wire xformtmp1639;
	assign xformtmp1639 = in[59] & in[743];
	wire xformtmp1589;
	assign xformtmp1589 = in[555] & xformtmp1639;
	wire xformtmp1380;
	assign xformtmp1380 = in[484] | xformtmp1589;
	wire xformtmp1551;
	assign xformtmp1551 = in[212] | xformtmp1380;
	wire xformtmp1733;
	assign xformtmp1733 = in[405] | xformtmp1551;
	wire xformtmp1832;
	assign xformtmp1832 = in[94] | in[940];
	wire xformtmp2068;
	assign xformtmp2068 = in[861] ^ xformtmp1832;
	wire xformtmp2162;
	assign xformtmp2162 = in[132] | xformtmp2068;
	wire xformtmp1518;
	assign xformtmp1518 = xformtmp1733 ^ xformtmp2162;
	wire xformtmp2146;
	assign xformtmp2146 = xformtmp1495 & xformtmp1518;
	wire xformtmp1461;
	assign xformtmp1461 = xformtmp1386 ^ xformtmp2146;
	wire xformtmp2248;
	assign xformtmp2248 = in[3] & in[175];
	wire xformtmp2105;
	assign xformtmp2105 = in[845] ^ xformtmp2248;
	wire xformtmp2234;
	assign xformtmp2234 = in[475] & xformtmp2105;
	wire xformtmp1296;
	assign xformtmp1296 = in[1151] ^ xformtmp2234;
	wire xformtmp1547;
	assign xformtmp1547 = in[835] | xformtmp1296;
	wire xformtmp1915;
	assign xformtmp1915 = in[111] ^ in[1284];
	wire xformtmp1501;
	assign xformtmp1501 = xformtmp1547 | xformtmp1915;
	wire xformtmp1674;
	assign xformtmp1674 = xformtmp1461 & xformtmp1501;
	wire xformtmp1981;
	assign xformtmp1981 = in[1086] & in[1214];
	wire xformtmp2171;
	assign xformtmp2171 = in[440] & xformtmp1981;
	wire xformtmp1646;
	assign xformtmp1646 = in[934] & xformtmp2171;
	wire xformtmp1758;
	assign xformtmp1758 = in[433] ^ in[745];
	wire xformtmp2093;
	assign xformtmp2093 = in[448] | in[641];
	wire xformtmp2218;
	assign xformtmp2218 = in[226] | xformtmp2093;
	wire xformtmp1895;
	assign xformtmp1895 = xformtmp1758 & xformtmp2218;
	wire xformtmp1976;
	assign xformtmp1976 = in[1071] ^ xformtmp1895;
	wire xformtmp1254;
	assign xformtmp1254 = xformtmp1646 ^ xformtmp1976;
	wire xformtmp1799;
	assign xformtmp1799 = in[174] ^ in[1232];
	wire xformtmp1911;
	assign xformtmp1911 = in[923] ^ xformtmp1799;
	wire xformtmp2168;
	assign xformtmp2168 = in[319] ^ in[924];
	wire xformtmp1692;
	assign xformtmp1692 = xformtmp1911 ^ xformtmp2168;
	wire xformtmp2187;
	assign xformtmp2187 = in[442] | xformtmp1692;
	wire xformtmp1643;
	assign xformtmp1643 = xformtmp1254 ^ xformtmp2187;
	wire xformtmp2195;
	assign xformtmp2195 = in[1199] ^ in[1245];
	wire xformtmp2063;
	assign xformtmp2063 = in[304] & in[586];
	wire xformtmp1853;
	assign xformtmp1853 = in[1231] | xformtmp2063;
	wire xformtmp1354;
	assign xformtmp1354 = in[187] | xformtmp1853;
	wire xformtmp1549;
	assign xformtmp1549 = in[26] ^ in[295];
	wire xformtmp1699;
	assign xformtmp1699 = xformtmp1354 & xformtmp1549;
	wire xformtmp1556;
	assign xformtmp1556 = in[84] | in[1119];
	wire xformtmp1985;
	assign xformtmp1985 = in[1017] ^ in[1326];
	wire xformtmp1859;
	assign xformtmp1859 = xformtmp1556 ^ xformtmp1985;
	wire xformtmp1303;
	assign xformtmp1303 = in[11] | xformtmp1859;
	wire xformtmp1878;
	assign xformtmp1878 = in[909] & in[918];
	wire xformtmp1936;
	assign xformtmp1936 = xformtmp1303 ^ xformtmp1878;
	wire xformtmp1512;
	assign xformtmp1512 = xformtmp1699 | xformtmp1936;
	wire xformtmp1836;
	assign xformtmp1836 = in[592] ^ in[937];
	wire xformtmp1817;
	assign xformtmp1817 = in[854] | xformtmp1836;
	wire xformtmp1640;
	assign xformtmp1640 = in[774] | in[1496];
	wire xformtmp2113;
	assign xformtmp2113 = in[819] ^ xformtmp1640;
	wire xformtmp1282;
	assign xformtmp1282 = xformtmp1817 | xformtmp2113;
	wire xformtmp1367;
	assign xformtmp1367 = in[167] | in[876];
	wire xformtmp2143;
	assign xformtmp2143 = in[1381] & xformtmp1367;
	wire xformtmp1457;
	assign xformtmp1457 = xformtmp1282 | xformtmp2143;
	wire xformtmp1898;
	assign xformtmp1898 = in[746] ^ in[1325];
	wire xformtmp2145;
	assign xformtmp2145 = xformtmp1457 | xformtmp1898;
	wire xformtmp1652;
	assign xformtmp1652 = xformtmp1512 & xformtmp2145;
	wire xformtmp1794;
	assign xformtmp1794 = in[45] ^ in[1261];
	wire xformtmp2198;
	assign xformtmp2198 = xformtmp1652 & xformtmp1794;
	wire xformtmp2156;
	assign xformtmp2156 = xformtmp2195 ^ xformtmp2198;
	wire xformtmp1888;
	assign xformtmp1888 = xformtmp1643 ^ xformtmp2156;
	wire xformtmp2124;
	assign xformtmp2124 = in[371] | in[1301];
	wire xformtmp1681;
	assign xformtmp1681 = in[666] ^ xformtmp2124;
	wire xformtmp1868;
	assign xformtmp1868 = in[1108] | xformtmp1681;
	wire xformtmp1595;
	assign xformtmp1595 = in[250] ^ xformtmp1868;
	wire xformtmp1789;
	assign xformtmp1789 = in[306] ^ in[623];
	wire xformtmp1931;
	assign xformtmp1931 = in[329] | xformtmp1789;
	wire xformtmp1466;
	assign xformtmp1466 = xformtmp1595 ^ xformtmp1931;
	wire xformtmp1345;
	assign xformtmp1345 = in[493] | xformtmp1466;
	wire xformtmp1416;
	assign xformtmp1416 = in[200] & in[855];
	wire xformtmp1920;
	assign xformtmp1920 = in[673] & in[1043];
	wire xformtmp1581;
	assign xformtmp1581 = in[253] ^ xformtmp1920;
	wire xformtmp1627;
	assign xformtmp1627 = in[675] ^ in[1260];
	wire xformtmp2131;
	assign xformtmp2131 = in[769] & xformtmp1627;
	wire xformtmp1352;
	assign xformtmp1352 = xformtmp1581 | xformtmp2131;
	wire xformtmp2225;
	assign xformtmp2225 = in[739] ^ in[791];
	wire xformtmp1815;
	assign xformtmp1815 = xformtmp1352 | xformtmp2225;
	wire xformtmp1667;
	assign xformtmp1667 = xformtmp1416 & xformtmp1815;
	wire xformtmp1948;
	assign xformtmp1948 = in[646] & xformtmp1667;
	wire xformtmp1329;
	assign xformtmp1329 = xformtmp1345 & xformtmp1948;
	wire xformtmp1500;
	assign xformtmp1500 = in[157] | in[974];
	wire xformtmp1972;
	assign xformtmp1972 = in[1285] | xformtmp1500;
	wire xformtmp1544;
	assign xformtmp1544 = in[594] & xformtmp1972;
	wire xformtmp2240;
	assign xformtmp2240 = in[50] & in[517];
	wire xformtmp1606;
	assign xformtmp1606 = in[788] ^ xformtmp2240;
	wire xformtmp2132;
	assign xformtmp2132 = xformtmp1544 & xformtmp1606;
	wire xformtmp1729;
	assign xformtmp1729 = in[234] ^ xformtmp2132;
	wire xformtmp2130;
	assign xformtmp2130 = in[929] & in[1483];
	wire xformtmp1749;
	assign xformtmp1749 = in[1493] ^ xformtmp2130;
	wire xformtmp1872;
	assign xformtmp1872 = in[408] & xformtmp1749;
	wire xformtmp1332;
	assign xformtmp1332 = xformtmp1729 ^ xformtmp1872;
	wire xformtmp2002;
	assign xformtmp2002 = xformtmp1329 ^ xformtmp1332;
	wire xformtmp2136;
	assign xformtmp2136 = xformtmp1888 | xformtmp2002;
	wire xformtmp1693;
	assign xformtmp1693 = in[824] ^ in[1083];
	wire xformtmp1423;
	assign xformtmp1423 = in[596] ^ in[996];
	wire xformtmp1866;
	assign xformtmp1866 = in[618] | in[1427];
	wire xformtmp1450;
	assign xformtmp1450 = in[450] & in[755];
	wire xformtmp2140;
	assign xformtmp2140 = in[215] | in[690];
	wire xformtmp2012;
	assign xformtmp2012 = in[438] & xformtmp2140;
	wire xformtmp1954;
	assign xformtmp1954 = xformtmp1450 & xformtmp2012;
	wire xformtmp2060;
	assign xformtmp2060 = xformtmp1866 | xformtmp1954;
	wire xformtmp1957;
	assign xformtmp1957 = xformtmp1423 | xformtmp2060;
	wire xformtmp1784;
	assign xformtmp1784 = in[1156] | xformtmp1957;
	wire xformtmp1481;
	assign xformtmp1481 = in[465] ^ xformtmp1784;
	wire xformtmp1801;
	assign xformtmp1801 = in[790] | in[1428];
	wire xformtmp1869;
	assign xformtmp1869 = in[783] & in[1080];
	wire xformtmp1827;
	assign xformtmp1827 = xformtmp1801 & xformtmp1869;
	wire xformtmp1427;
	assign xformtmp1427 = in[655] | xformtmp1827;
	wire xformtmp1656;
	assign xformtmp1656 = in[292] | xformtmp1427;
	wire xformtmp1945;
	assign xformtmp1945 = xformtmp1481 | xformtmp1656;
	wire xformtmp1256;
	assign xformtmp1256 = in[238] & in[1476];
	wire xformtmp1995;
	assign xformtmp1995 = in[773] ^ xformtmp1256;
	wire xformtmp1609;
	assign xformtmp1609 = xformtmp1945 ^ xformtmp1995;
	wire xformtmp2005;
	assign xformtmp2005 = in[722] ^ xformtmp1609;
	wire xformtmp1558;
	assign xformtmp1558 = xformtmp1693 & xformtmp2005;
	wire xformtmp1394;
	assign xformtmp1394 = in[6] ^ in[629];
	wire xformtmp1339;
	assign xformtmp1339 = in[1452] & xformtmp1394;
	wire xformtmp2008;
	assign xformtmp2008 = in[219] & xformtmp1339;
	wire xformtmp1486;
	assign xformtmp1486 = in[54] & xformtmp2008;
	wire xformtmp1276;
	assign xformtmp1276 = in[568] & in[1442];
	wire xformtmp1534;
	assign xformtmp1534 = in[689] & xformtmp1276;
	wire xformtmp1519;
	assign xformtmp1519 = in[1235] & in[1389];
	wire xformtmp1992;
	assign xformtmp1992 = in[181] | xformtmp1519;
	wire xformtmp1765;
	assign xformtmp1765 = xformtmp1534 ^ xformtmp1992;
	wire xformtmp1642;
	assign xformtmp1642 = xformtmp1486 ^ xformtmp1765;
	wire xformtmp2201;
	assign xformtmp2201 = in[86] | in[407];
	wire xformtmp1763;
	assign xformtmp1763 = in[103] & xformtmp2201;
	wire xformtmp2029;
	assign xformtmp2029 = in[291] ^ in[705];
	wire xformtmp1881;
	assign xformtmp1881 = in[125] & xformtmp2029;
	wire xformtmp1564;
	assign xformtmp1564 = xformtmp1763 ^ xformtmp1881;
	wire xformtmp1741;
	assign xformtmp1741 = in[107] | in[740];
	wire xformtmp1964;
	assign xformtmp1964 = in[1054] & xformtmp1741;
	wire xformtmp1585;
	assign xformtmp1585 = xformtmp1564 | xformtmp1964;
	wire xformtmp2016;
	assign xformtmp2016 = in[302] ^ in[1148];
	wire xformtmp1304;
	assign xformtmp1304 = in[1144] & xformtmp2016;
	wire xformtmp1766;
	assign xformtmp1766 = in[648] | in[1449];
	wire xformtmp1406;
	assign xformtmp1406 = in[619] ^ xformtmp1766;
	wire xformtmp1850;
	assign xformtmp1850 = xformtmp1304 & xformtmp1406;
	wire xformtmp1909;
	assign xformtmp1909 = in[723] | in[821];
	wire xformtmp1648;
	assign xformtmp1648 = xformtmp1850 | xformtmp1909;
	wire xformtmp1730;
	assign xformtmp1730 = in[161] | in[1166];
	wire xformtmp1307;
	assign xformtmp1307 = in[864] ^ xformtmp1730;
	wire xformtmp2116;
	assign xformtmp2116 = in[404] ^ in[1130];
	wire xformtmp2137;
	assign xformtmp2137 = in[145] ^ in[299];
	wire xformtmp1550;
	assign xformtmp1550 = xformtmp2116 ^ xformtmp2137;
	wire xformtmp2014;
	assign xformtmp2014 = in[349] ^ in[1307];
	wire xformtmp1616;
	assign xformtmp1616 = in[778] ^ xformtmp2014;
	wire xformtmp2249;
	assign xformtmp2249 = xformtmp1550 & xformtmp1616;
	wire xformtmp1852;
	assign xformtmp1852 = xformtmp1307 & xformtmp2249;
	wire xformtmp1588;
	assign xformtmp1588 = in[73] & in[1327];
	wire xformtmp1917;
	assign xformtmp1917 = in[1195] & xformtmp1588;
	wire xformtmp2233;
	assign xformtmp2233 = in[1135] & xformtmp1917;
	wire xformtmp1715;
	assign xformtmp1715 = xformtmp1852 & xformtmp2233;
	wire xformtmp1778;
	assign xformtmp1778 = xformtmp1648 ^ xformtmp1715;
	wire xformtmp1502;
	assign xformtmp1502 = in[92] & xformtmp1778;
	wire xformtmp1891;
	assign xformtmp1891 = in[1027] | in[1177];
	wire xformtmp2114;
	assign xformtmp2114 = in[730] & xformtmp1891;
	wire xformtmp2191;
	assign xformtmp2191 = in[1057] | xformtmp2114;
	wire xformtmp1487;
	assign xformtmp1487 = in[1154] & xformtmp2191;
	wire xformtmp2206;
	assign xformtmp2206 = in[476] ^ xformtmp1487;
	wire xformtmp1448;
	assign xformtmp1448 = xformtmp1502 ^ xformtmp2206;
	wire xformtmp1701;
	assign xformtmp1701 = in[1041] | in[1306];
	wire xformtmp1513;
	assign xformtmp1513 = in[118] & in[1182];
	wire xformtmp1792;
	assign xformtmp1792 = in[563] ^ xformtmp1513;
	wire xformtmp1880;
	assign xformtmp1880 = in[1407] | xformtmp1792;
	wire xformtmp1727;
	assign xformtmp1727 = xformtmp1701 | xformtmp1880;
	wire xformtmp1664;
	assign xformtmp1664 = xformtmp1448 ^ xformtmp1727;
	wire xformtmp1465;
	assign xformtmp1465 = xformtmp1585 ^ xformtmp1664;
	wire xformtmp1533;
	assign xformtmp1533 = in[803] ^ in[1175];
	wire xformtmp1634;
	assign xformtmp1634 = in[954] ^ xformtmp1533;
	wire xformtmp2056;
	assign xformtmp2056 = in[80] & in[284];
	wire xformtmp1822;
	assign xformtmp1822 = in[471] ^ xformtmp2056;
	wire xformtmp1433;
	assign xformtmp1433 = xformtmp1634 ^ xformtmp1822;
	wire xformtmp1372;
	assign xformtmp1372 = in[179] ^ in[753];
	wire xformtmp1462;
	assign xformtmp1462 = in[246] & xformtmp1372;
	wire xformtmp1777;
	assign xformtmp1777 = in[385] & in[1349];
	wire xformtmp2039;
	assign xformtmp2039 = in[865] | in[1058];
	wire xformtmp2237;
	assign xformtmp2237 = in[889] ^ xformtmp2039;
	wire xformtmp1918;
	assign xformtmp1918 = in[603] & xformtmp2237;
	wire xformtmp1828;
	assign xformtmp1828 = xformtmp1777 ^ xformtmp1918;
	wire xformtmp1243;
	assign xformtmp1243 = xformtmp1462 | xformtmp1828;
	wire xformtmp1374;
	assign xformtmp1374 = in[528] & in[1112];
	wire xformtmp1900;
	assign xformtmp1900 = in[490] ^ xformtmp1374;
	wire xformtmp1514;
	assign xformtmp1514 = in[1487] & xformtmp1900;
	wire xformtmp1568;
	assign xformtmp1568 = in[216] | in[419];
	wire xformtmp1604;
	assign xformtmp1604 = in[1287] ^ xformtmp1568;
	wire xformtmp1944;
	assign xformtmp1944 = in[268] ^ xformtmp1604;
	wire xformtmp1764;
	assign xformtmp1764 = in[1001] & xformtmp1944;
	wire xformtmp1607;
	assign xformtmp1607 = xformtmp1514 | xformtmp1764;
	wire xformtmp1522;
	assign xformtmp1522 = in[1422] ^ xformtmp1607;
	wire xformtmp1965;
	assign xformtmp1965 = xformtmp1243 & xformtmp1522;
	wire xformtmp1759;
	assign xformtmp1759 = xformtmp1433 & xformtmp1965;
	wire xformtmp1317;
	assign xformtmp1317 = xformtmp1465 ^ xformtmp1759;
	wire xformtmp1503;
	assign xformtmp1503 = in[968] | in[1418];
	wire xformtmp2106;
	assign xformtmp2106 = in[998] & xformtmp1503;
	wire xformtmp2239;
	assign xformtmp2239 = in[142] & in[919];
	wire xformtmp1983;
	assign xformtmp1983 = xformtmp2106 ^ xformtmp2239;
	wire xformtmp2030;
	assign xformtmp2030 = in[1340] | xformtmp1983;
	wire xformtmp2072;
	assign xformtmp2072 = in[887] & xformtmp2030;
	wire xformtmp1717;
	assign xformtmp1717 = xformtmp1317 | xformtmp2072;
	wire xformtmp1548;
	assign xformtmp1548 = xformtmp1642 ^ xformtmp1717;
	wire xformtmp1483;
	assign xformtmp1483 = in[261] | in[324];
	wire xformtmp1520;
	assign xformtmp1520 = in[195] & in[570];
	wire xformtmp1497;
	assign xformtmp1497 = in[467] ^ xformtmp1520;
	wire xformtmp1835;
	assign xformtmp1835 = in[69] & in[355];
	wire xformtmp1795;
	assign xformtmp1795 = xformtmp1497 | xformtmp1835;
	wire xformtmp2220;
	assign xformtmp2220 = xformtmp1483 & xformtmp1795;
	wire xformtmp2251;
	assign xformtmp2251 = xformtmp1548 ^ xformtmp2220;
	wire xformtmp2256;
	assign xformtmp2256 = xformtmp1558 | xformtmp2251;
	wire xformtmp1816;
	assign xformtmp1816 = xformtmp2136 & xformtmp2256;
	wire xformtmp1578;
	assign xformtmp1578 = xformtmp1674 | xformtmp1816;
	wire xformtmp2051;
	assign xformtmp2051 = in[1376] ^ in[1473];
	wire xformtmp1553;
	assign xformtmp1553 = in[1457] | xformtmp2051;
	wire xformtmp1400;
	assign xformtmp1400 = in[336] | in[579];
	wire xformtmp1454;
	assign xformtmp1454 = in[267] ^ in[1242];
	wire xformtmp1724;
	assign xformtmp1724 = in[469] & in[573];
	wire xformtmp1747;
	assign xformtmp1747 = xformtmp1454 | xformtmp1724;
	wire xformtmp1555;
	assign xformtmp1555 = xformtmp1400 & xformtmp1747;
	wire xformtmp1479;
	assign xformtmp1479 = in[141] & xformtmp1555;
	wire xformtmp1812;
	assign xformtmp1812 = in[113] ^ in[958];
	wire xformtmp1949;
	assign xformtmp1949 = xformtmp1479 | xformtmp1812;
	wire xformtmp1405;
	assign xformtmp1405 = xformtmp1553 & xformtmp1949;
	wire xformtmp1444;
	assign xformtmp1444 = in[296] ^ in[1303];
	wire xformtmp1618;
	assign xformtmp1618 = in[844] ^ xformtmp1444;
	wire xformtmp1521;
	assign xformtmp1521 = xformtmp1405 ^ xformtmp1618;
	wire xformtmp1273;
	assign xformtmp1273 = in[49] ^ in[713];
	wire xformtmp1244;
	assign xformtmp1244 = in[1059] ^ in[1075];
	wire xformtmp1603;
	assign xformtmp1603 = in[1341] ^ in[1406];
	wire xformtmp2038;
	assign xformtmp2038 = in[699] | in[1040];
	wire xformtmp2111;
	assign xformtmp2111 = xformtmp1603 | xformtmp2038;
	wire xformtmp2058;
	assign xformtmp2058 = xformtmp1244 | xformtmp2111;
	wire xformtmp1403;
	assign xformtmp1403 = xformtmp1273 ^ xformtmp2058;
	wire xformtmp1608;
	assign xformtmp1608 = in[925] ^ xformtmp1403;
	wire xformtmp1531;
	assign xformtmp1531 = in[1443] ^ xformtmp1608;
	wire xformtmp2188;
	assign xformtmp2188 = in[283] ^ xformtmp1531;
	wire xformtmp1601;
	assign xformtmp1601 = xformtmp1521 ^ xformtmp2188;
	wire xformtmp1325;
	assign xformtmp1325 = in[485] & in[1159];
	wire xformtmp2065;
	assign xformtmp2065 = in[1023] ^ in[1342];
	wire xformtmp1541;
	assign xformtmp1541 = in[969] ^ xformtmp2065;
	wire xformtmp1395;
	assign xformtmp1395 = in[1425] | xformtmp1541;
	wire xformtmp1813;
	assign xformtmp1813 = xformtmp1325 & xformtmp1395;
	wire xformtmp1562;
	assign xformtmp1562 = in[39] & xformtmp1813;
	wire xformtmp1341;
	assign xformtmp1341 = in[260] | in[1267];
	wire xformtmp2094;
	assign xformtmp2094 = in[637] | in[826];
	wire xformtmp1343;
	assign xformtmp1343 = xformtmp1341 ^ xformtmp2094;
	wire xformtmp2032;
	assign xformtmp2032 = in[994] | in[1365];
	wire xformtmp1290;
	assign xformtmp1290 = xformtmp1343 & xformtmp2032;
	wire xformtmp1418;
	assign xformtmp1418 = in[1420] & in[1430];
	wire xformtmp2215;
	assign xformtmp2215 = xformtmp1290 ^ xformtmp1418;
	wire xformtmp1583;
	assign xformtmp1583 = in[352] ^ xformtmp2215;
	wire xformtmp1361;
	assign xformtmp1361 = xformtmp1562 | xformtmp1583;
	wire xformtmp2047;
	assign xformtmp2047 = in[667] & in[793];
	wire xformtmp1809;
	assign xformtmp1809 = in[483] | xformtmp2047;
	wire xformtmp1847;
	assign xformtmp1847 = in[616] | xformtmp1809;
	wire xformtmp1314;
	assign xformtmp1314 = in[43] ^ xformtmp1847;
	wire xformtmp1984;
	assign xformtmp1984 = in[552] | in[1046];
	wire xformtmp2189;
	assign xformtmp2189 = in[147] ^ xformtmp1984;
	wire xformtmp1382;
	assign xformtmp1382 = xformtmp1314 ^ xformtmp2189;
	wire xformtmp1302;
	assign xformtmp1302 = in[1405] ^ xformtmp1382;
	wire xformtmp2226;
	assign xformtmp2226 = in[198] & in[588];
	wire xformtmp1360;
	assign xformtmp1360 = in[693] & xformtmp2226;
	wire xformtmp1348;
	assign xformtmp1348 = in[25] ^ xformtmp1360;
	wire xformtmp1572;
	assign xformtmp1572 = in[1481] | xformtmp1348;
	wire xformtmp1288;
	assign xformtmp1288 = in[75] & xformtmp1572;
	wire xformtmp1873;
	assign xformtmp1873 = in[515] | in[1468];
	wire xformtmp1644;
	assign xformtmp1644 = xformtmp1288 ^ xformtmp1873;
	wire xformtmp1744;
	assign xformtmp1744 = in[565] | in[1308];
	wire xformtmp1245;
	assign xformtmp1245 = in[744] ^ xformtmp1744;
	wire xformtmp1459;
	assign xformtmp1459 = in[587] ^ xformtmp1245;
	wire xformtmp1399;
	assign xformtmp1399 = in[71] & in[192];
	wire xformtmp1933;
	assign xformtmp1933 = in[967] ^ xformtmp1399;
	wire xformtmp1754;
	assign xformtmp1754 = in[236] ^ in[1181];
	wire xformtmp1482;
	assign xformtmp1482 = in[1391] ^ xformtmp1754;
	wire xformtmp2035;
	assign xformtmp2035 = in[1076] & xformtmp1482;
	wire xformtmp1829;
	assign xformtmp1829 = xformtmp1933 ^ xformtmp2035;
	wire xformtmp2244;
	assign xformtmp2244 = in[290] ^ in[1374];
	wire xformtmp1688;
	assign xformtmp1688 = in[684] & xformtmp2244;
	wire xformtmp2151;
	assign xformtmp2151 = in[1290] | xformtmp1688;
	wire xformtmp1308;
	assign xformtmp1308 = xformtmp1829 & xformtmp2151;
	wire xformtmp2083;
	assign xformtmp2083 = in[1078] | in[1388];
	wire xformtmp2184;
	assign xformtmp2184 = in[140] ^ in[1484];
	wire xformtmp1732;
	assign xformtmp1732 = xformtmp2083 & xformtmp2184;
	wire xformtmp1980;
	assign xformtmp1980 = in[16] | xformtmp1732;
	wire xformtmp1437;
	assign xformtmp1437 = in[254] ^ in[487];
	wire xformtmp2169;
	assign xformtmp2169 = in[893] & xformtmp1437;
	wire xformtmp1756;
	assign xformtmp1756 = xformtmp1980 ^ xformtmp2169;
	wire xformtmp1358;
	assign xformtmp1358 = xformtmp1308 & xformtmp1756;
	wire xformtmp1430;
	assign xformtmp1430 = in[170] ^ in[736];
	wire xformtmp1364;
	assign xformtmp1364 = in[323] | in[858];
	wire xformtmp1755;
	assign xformtmp1755 = in[205] | in[547];
	wire xformtmp1772;
	assign xformtmp1772 = xformtmp1364 | xformtmp1755;
	wire xformtmp2073;
	assign xformtmp2073 = xformtmp1430 | xformtmp1772;
	wire xformtmp2242;
	assign xformtmp2242 = xformtmp1358 ^ xformtmp2073;
	wire xformtmp2250;
	assign xformtmp2250 = xformtmp1459 & xformtmp2242;
	wire xformtmp1857;
	assign xformtmp1857 = xformtmp1644 | xformtmp2250;
	wire xformtmp1671;
	assign xformtmp1671 = xformtmp1302 | xformtmp1857;
	wire xformtmp1428;
	assign xformtmp1428 = in[325] | in[1184];
	wire xformtmp1523;
	assign xformtmp1523 = in[696] & xformtmp1428;
	wire xformtmp1855;
	assign xformtmp1855 = in[712] & xformtmp1523;
	wire xformtmp1804;
	assign xformtmp1804 = in[559] | xformtmp1855;
	wire xformtmp1480;
	assign xformtmp1480 = xformtmp1671 | xformtmp1804;
	wire xformtmp1951;
	assign xformtmp1951 = xformtmp1361 ^ xformtmp1480;
	wire xformtmp1922;
	assign xformtmp1922 = xformtmp1601 | xformtmp1951;
	wire xformtmp2235;
	assign xformtmp2235 = xformtmp1578 | xformtmp1922;
	wire xformtmp1439;
	assign xformtmp1439 = xformtmp1660 ^ xformtmp2235;
	wire xformtmp1280;
	assign xformtmp1280 = in[1283] & in[1375];
	wire xformtmp1808;
	assign xformtmp1808 = in[204] | in[532];
	wire xformtmp1958;
	assign xformtmp1958 = in[1321] & xformtmp1808;
	wire xformtmp1926;
	assign xformtmp1926 = in[1068] ^ in[1410];
	wire xformtmp1326;
	assign xformtmp1326 = in[698] ^ xformtmp1926;
	wire xformtmp1426;
	assign xformtmp1426 = in[121] | in[1125];
	wire xformtmp1613;
	assign xformtmp1613 = in[308] & xformtmp1426;
	wire xformtmp1978;
	assign xformtmp1978 = in[1469] & xformtmp1613;
	wire xformtmp2160;
	assign xformtmp2160 = xformtmp1326 ^ xformtmp1978;
	wire xformtmp2170;
	assign xformtmp2170 = xformtmp1958 | xformtmp2160;
	wire xformtmp1499;
	assign xformtmp1499 = in[88] | in[1482];
	wire xformtmp2112;
	assign xformtmp2112 = in[287] ^ xformtmp1499;
	wire xformtmp1890;
	assign xformtmp1890 = in[1330] & xformtmp2112;
	wire xformtmp1552;
	assign xformtmp1552 = in[683] & in[732];
	wire xformtmp2097;
	assign xformtmp2097 = in[657] ^ in[801];
	wire xformtmp2219;
	assign xformtmp2219 = xformtmp1552 ^ xformtmp2097;
	wire xformtmp1679;
	assign xformtmp1679 = xformtmp1890 ^ xformtmp2219;
	wire xformtmp1737;
	assign xformtmp1737 = in[578] | in[1455];
	wire xformtmp1824;
	assign xformtmp1824 = in[1219] ^ xformtmp1737;
	wire xformtmp2217;
	assign xformtmp2217 = xformtmp1679 ^ xformtmp1824;
	wire xformtmp1826;
	assign xformtmp1826 = xformtmp2170 ^ xformtmp2217;
	wire xformtmp1956;
	assign xformtmp1956 = in[1282] & in[1288];
	wire xformtmp1241;
	assign xformtmp1241 = in[343] | in[711];
	wire xformtmp2243;
	assign xformtmp2243 = in[37] | in[1431];
	wire xformtmp2148;
	assign xformtmp2148 = xformtmp1241 & xformtmp2243;
	wire xformtmp2221;
	assign xformtmp2221 = in[668] & in[1390];
	wire xformtmp2055;
	assign xformtmp2055 = xformtmp2148 & xformtmp2221;
	wire xformtmp1901;
	assign xformtmp1901 = xformtmp1956 ^ xformtmp2055;
	wire xformtmp1347;
	assign xformtmp1347 = in[351] & in[674];
	wire xformtmp1388;
	assign xformtmp1388 = in[1085] & xformtmp1347;
	wire xformtmp2121;
	assign xformtmp2121 = in[700] ^ in[1176];
	wire xformtmp2133;
	assign xformtmp2133 = xformtmp1388 ^ xformtmp2121;
	wire xformtmp2134;
	assign xformtmp2134 = in[1066] ^ in[1070];
	wire xformtmp2082;
	assign xformtmp2082 = xformtmp2133 ^ xformtmp2134;
	wire xformtmp1979;
	assign xformtmp1979 = xformtmp1901 & xformtmp2082;
	wire xformtmp2075;
	assign xformtmp2075 = xformtmp1826 ^ xformtmp1979;
	wire xformtmp1821;
	assign xformtmp1821 = xformtmp1280 | xformtmp2075;
	wire xformtmp1258;
	assign xformtmp1258 = in[232] | in[1222];
	wire xformtmp1536;
	assign xformtmp1536 = in[337] | in[1049];
	wire xformtmp1990;
	assign xformtmp1990 = xformtmp1258 & xformtmp1536;
	wire xformtmp1340;
	assign xformtmp1340 = in[1165] & in[1189];
	wire xformtmp2026;
	assign xformtmp2026 = in[1396] ^ xformtmp1340;
	wire xformtmp1787;
	assign xformtmp1787 = in[678] ^ in[1300];
	wire xformtmp2031;
	assign xformtmp2031 = in[540] | xformtmp1787;
	wire xformtmp1508;
	assign xformtmp1508 = xformtmp2026 | xformtmp2031;
	wire xformtmp1420;
	assign xformtmp1420 = in[190] & in[449];
	wire xformtmp1968;
	assign xformtmp1968 = in[617] & in[880];
	wire xformtmp1617;
	assign xformtmp1617 = xformtmp1420 | xformtmp1968;
	wire xformtmp2087;
	assign xformtmp2087 = xformtmp1508 | xformtmp1617;
	wire xformtmp1493;
	assign xformtmp1493 = xformtmp1990 & xformtmp2087;
	wire xformtmp1938;
	assign xformtmp1938 = in[416] | in[1262];
	wire xformtmp1955;
	assign xformtmp1955 = xformtmp1493 & xformtmp1938;
	wire xformtmp2034;
	assign xformtmp2034 = in[100] | in[1343];
	wire xformtmp2127;
	assign xformtmp2127 = in[272] & in[435];
	wire xformtmp2099;
	assign xformtmp2099 = xformtmp2034 | xformtmp2127;
	wire xformtmp1914;
	assign xformtmp1914 = in[395] & in[656];
	wire xformtmp1344;
	assign xformtmp1344 = in[393] | xformtmp1914;
	wire xformtmp1840;
	assign xformtmp1840 = in[311] | xformtmp1344;
	wire xformtmp2049;
	assign xformtmp2049 = in[109] ^ in[805];
	wire xformtmp2149;
	assign xformtmp2149 = xformtmp1840 | xformtmp2049;
	wire xformtmp1526;
	assign xformtmp1526 = xformtmp2099 | xformtmp2149;
	wire xformtmp1662;
	assign xformtmp1662 = in[184] & in[259];
	wire xformtmp1369;
	assign xformtmp1369 = in[307] & in[1221];
	wire xformtmp1742;
	assign xformtmp1742 = in[1019] | in[1185];
	wire xformtmp2023;
	assign xformtmp2023 = xformtmp1369 ^ xformtmp1742;
	wire xformtmp1993;
	assign xformtmp1993 = in[277] ^ xformtmp2023;
	wire xformtmp2181;
	assign xformtmp2181 = in[415] | in[1011];
	wire xformtmp1885;
	assign xformtmp1885 = xformtmp1993 & xformtmp2181;
	wire xformtmp1464;
	assign xformtmp1464 = in[178] & in[871];
	wire xformtmp1728;
	assign xformtmp1728 = in[497] | in[1088];
	wire xformtmp1540;
	assign xformtmp1540 = in[60] | xformtmp1728;
	wire xformtmp1424;
	assign xformtmp1424 = xformtmp1464 & xformtmp1540;
	wire xformtmp2199;
	assign xformtmp2199 = in[76] & in[622];
	wire xformtmp1930;
	assign xformtmp1930 = xformtmp1424 | xformtmp2199;
	wire xformtmp1823;
	assign xformtmp1823 = xformtmp1885 ^ xformtmp1930;
	wire xformtmp1292;
	assign xformtmp1292 = in[965] | xformtmp1823;
	wire xformtmp1381;
	assign xformtmp1381 = in[499] | in[527];
	wire xformtmp1496;
	assign xformtmp1496 = xformtmp1292 | xformtmp1381;
	wire xformtmp1321;
	assign xformtmp1321 = in[556] & in[1079];
	wire xformtmp1271;
	assign xformtmp1271 = in[144] | xformtmp1321;
	wire xformtmp2119;
	assign xformtmp2119 = in[526] ^ xformtmp1271;
	wire xformtmp1431;
	assign xformtmp1431 = in[859] ^ xformtmp2119;
	wire xformtmp1861;
	assign xformtmp1861 = in[945] | in[975];
	wire xformtmp2045;
	assign xformtmp2045 = xformtmp1431 ^ xformtmp1861;
	wire xformtmp1327;
	assign xformtmp1327 = xformtmp1496 | xformtmp2045;
	wire xformtmp1743;
	assign xformtmp1743 = in[888] | in[1352];
	wire xformtmp1769;
	assign xformtmp1769 = in[849] & in[1461];
	wire xformtmp2017;
	assign xformtmp2017 = in[155] & in[671];
	wire xformtmp1894;
	assign xformtmp1894 = xformtmp1769 & xformtmp2017;
	wire xformtmp1260;
	assign xformtmp1260 = xformtmp1743 | xformtmp1894;
	wire xformtmp1690;
	assign xformtmp1690 = in[1163] | xformtmp1260;
	wire xformtmp2128;
	assign xformtmp2128 = xformtmp1327 ^ xformtmp1690;
	wire xformtmp1994;
	assign xformtmp1994 = xformtmp1662 ^ xformtmp2128;
	wire xformtmp2019;
	assign xformtmp2019 = xformtmp1526 ^ xformtmp1994;
	wire xformtmp1761;
	assign xformtmp1761 = xformtmp1955 & xformtmp2019;
	wire xformtmp2223;
	assign xformtmp2223 = in[1448] & in[1459];
	wire xformtmp1529;
	assign xformtmp1529 = xformtmp1761 & xformtmp2223;
	wire xformtmp2126;
	assign xformtmp2126 = in[249] ^ in[548];
	wire xformtmp1790;
	assign xformtmp1790 = in[85] & xformtmp2126;
	wire xformtmp1263;
	assign xformtmp1263 = in[806] & xformtmp1790;
	wire xformtmp1490;
	assign xformtmp1490 = in[218] ^ in[1358];
	wire xformtmp1262;
	assign xformtmp1262 = in[1265] | xformtmp1490;
	wire xformtmp1714;
	assign xformtmp1714 = in[67] & in[916];
	wire xformtmp1537;
	assign xformtmp1537 = in[309] & xformtmp1714;
	wire xformtmp1334;
	assign xformtmp1334 = xformtmp1262 | xformtmp1537;
	wire xformtmp1726;
	assign xformtmp1726 = in[42] & in[1370];
	wire xformtmp1469;
	assign xformtmp1469 = in[128] ^ xformtmp1726;
	wire xformtmp1443;
	assign xformtmp1443 = in[950] & xformtmp1469;
	wire xformtmp2080;
	assign xformtmp2080 = in[27] ^ in[437];
	wire xformtmp2154;
	assign xformtmp2154 = in[1279] & xformtmp2080;
	wire xformtmp1919;
	assign xformtmp1919 = xformtmp1443 | xformtmp2154;
	wire xformtmp1266;
	assign xformtmp1266 = xformtmp1334 & xformtmp1919;
	wire xformtmp1316;
	assign xformtmp1316 = xformtmp1263 | xformtmp1266;
	wire xformtmp1622;
	assign xformtmp1622 = in[30] & xformtmp1316;
	wire xformtmp1860;
	assign xformtmp1860 = in[608] & in[908];
	wire xformtmp1470;
	assign xformtmp1470 = in[134] & in[863];
	wire xformtmp1879;
	assign xformtmp1879 = in[538] & in[1359];
	wire xformtmp2074;
	assign xformtmp2074 = xformtmp1470 | xformtmp1879;
	wire xformtmp1867;
	assign xformtmp1867 = in[359] | xformtmp2074;
	wire xformtmp1401;
	assign xformtmp1401 = xformtmp1860 & xformtmp1867;
	wire xformtmp2091;
	assign xformtmp2091 = in[14] & in[638];
	wire xformtmp2053;
	assign xformtmp2053 = in[939] ^ xformtmp2091;
	wire xformtmp2152;
	assign xformtmp2152 = in[78] | xformtmp2053;
	wire xformtmp1543;
	assign xformtmp1543 = in[1116] ^ xformtmp2152;
	wire xformtmp1839;
	assign xformtmp1839 = in[19] | in[421];
	wire xformtmp2144;
	assign xformtmp2144 = in[628] ^ xformtmp1839;
	wire xformtmp1830;
	assign xformtmp1830 = in[1113] & xformtmp2144;
	wire xformtmp2007;
	assign xformtmp2007 = xformtmp1543 | xformtmp1830;
	wire xformtmp1731;
	assign xformtmp1731 = in[566] ^ xformtmp2007;
	wire xformtmp2129;
	assign xformtmp2129 = xformtmp1401 | xformtmp1731;
	wire xformtmp1745;
	assign xformtmp1745 = xformtmp1622 | xformtmp2129;
	wire xformtmp2102;
	assign xformtmp2102 = xformtmp1529 | xformtmp1745;
	wire xformtmp1905;
	assign xformtmp1905 = xformtmp1821 & xformtmp2102;
	wire xformtmp1471;
	assign xformtmp1471 = xformtmp1439 ^ xformtmp1905;
	wire xformtmp1474;
	assign xformtmp1474 = in[102] | in[664];
	wire xformtmp1781;
	assign xformtmp1781 = in[1247] ^ xformtmp1474;
	wire xformtmp1286;
	assign xformtmp1286 = in[577] | in[1441];
	wire xformtmp1532;
	assign xformtmp1532 = in[951] & xformtmp1286;
	wire xformtmp1338;
	assign xformtmp1338 = in[1150] ^ xformtmp1532;
	wire xformtmp2009;
	assign xformtmp2009 = in[305] | in[1180];
	wire xformtmp1982;
	assign xformtmp1982 = in[1146] ^ xformtmp2009;
	wire xformtmp1935;
	assign xformtmp1935 = in[1319] ^ xformtmp1982;
	wire xformtmp1863;
	assign xformtmp1863 = xformtmp1338 | xformtmp1935;
	wire xformtmp1963;
	assign xformtmp1963 = in[1356] | xformtmp1863;
	wire xformtmp1600;
	assign xformtmp1600 = xformtmp1781 & xformtmp1963;
	wire xformtmp1767;
	assign xformtmp1767 = in[32] & in[550];
	wire xformtmp1287;
	assign xformtmp1287 = xformtmp1600 & xformtmp1767;
	wire xformtmp1255;
	assign xformtmp1255 = in[902] | in[1280];
	wire xformtmp1579;
	assign xformtmp1579 = in[1432] | xformtmp1255;
	wire xformtmp1385;
	assign xformtmp1385 = in[1421] ^ xformtmp1579;
	wire xformtmp2166;
	assign xformtmp2166 = in[46] & in[333];
	wire xformtmp2098;
	assign xformtmp2098 = xformtmp1385 | xformtmp2166;
	wire xformtmp1686;
	assign xformtmp1686 = in[895] | in[1318];
	wire xformtmp1398;
	assign xformtmp1398 = in[143] ^ in[1200];
	wire xformtmp2037;
	assign xformtmp2037 = in[17] | xformtmp1398;
	wire xformtmp1842;
	assign xformtmp1842 = in[727] & xformtmp2037;
	wire xformtmp1434;
	assign xformtmp1434 = in[18] | xformtmp1842;
	wire xformtmp1837;
	assign xformtmp1837 = in[979] ^ xformtmp1434;
	wire xformtmp2107;
	assign xformtmp2107 = xformtmp1686 | xformtmp1837;
	wire xformtmp1599;
	assign xformtmp1599 = xformtmp2098 | xformtmp2107;
	wire xformtmp1377;
	assign xformtmp1377 = xformtmp1287 & xformtmp1599;
	wire xformtmp1333;
	assign xformtmp1333 = in[1009] & in[1128];
	wire xformtmp1940;
	assign xformtmp1940 = in[1031] ^ in[1351];
	wire xformtmp2042;
	assign xformtmp2042 = in[572] & xformtmp1940;
	wire xformtmp1899;
	assign xformtmp1899 = xformtmp1333 ^ xformtmp2042;
	wire xformtmp1267;
	assign xformtmp1267 = in[264] | xformtmp1899;
	wire xformtmp1638;
	assign xformtmp1638 = in[782] ^ in[878];
	wire xformtmp1557;
	assign xformtmp1557 = xformtmp1267 & xformtmp1638;
	wire xformtmp1586;
	assign xformtmp1586 = in[839] & in[1392];
	wire xformtmp2216;
	assign xformtmp2216 = in[262] & xformtmp1586;
	wire xformtmp1353;
	assign xformtmp1353 = in[453] | xformtmp2216;
	wire xformtmp1637;
	assign xformtmp1637 = in[798] ^ in[962];
	wire xformtmp2230;
	assign xformtmp2230 = xformtmp1353 & xformtmp1637;
	wire xformtmp1320;
	assign xformtmp1320 = xformtmp1557 ^ xformtmp2230;
	wire xformtmp1807;
	assign xformtmp1807 = in[424] ^ in[987];
	wire xformtmp2203;
	assign xformtmp2203 = in[663] & xformtmp1807;
	wire xformtmp1577;
	assign xformtmp1577 = in[418] | xformtmp2203;
	wire xformtmp1939;
	assign xformtmp1939 = in[1445] | xformtmp1577;
	wire xformtmp1628;
	assign xformtmp1628 = in[523] ^ in[1012];
	wire xformtmp2173;
	assign xformtmp2173 = in[1149] & xformtmp1628;
	wire xformtmp2178;
	assign xformtmp2178 = xformtmp1939 | xformtmp2173;
	wire xformtmp2163;
	assign xformtmp2163 = in[1162] & xformtmp2178;
	wire xformtmp2246;
	assign xformtmp2246 = xformtmp1320 | xformtmp2163;
	wire xformtmp1666;
	assign xformtmp1666 = xformtmp1377 ^ xformtmp2246;
	wire xformtmp1584;
	assign xformtmp1584 = xformtmp1471 | xformtmp1666;
	wire xformtmp1986;
	assign xformtmp1986 = xformtmp1441 ^ xformtmp1584;
	wire xformtmp1391;
	assign xformtmp1391 = xformtmp1538 & xformtmp1986;
	wire xformtmp1580;
	assign xformtmp1580 = in[61] & in[688];
	wire xformtmp1780;
	assign xformtmp1780 = in[964] ^ xformtmp1580;
	wire xformtmp1746;
	assign xformtmp1746 = in[1206] ^ xformtmp1780;
	wire xformtmp1750;
	assign xformtmp1750 = in[506] & xformtmp1746;
	wire xformtmp1912;
	assign xformtmp1912 = in[1207] & in[1354];
	wire xformtmp2081;
	assign xformtmp2081 = xformtmp1750 | xformtmp1912;
	wire xformtmp1265;
	assign xformtmp1265 = in[1337] ^ xformtmp2081;
	wire xformtmp1494;
	assign xformtmp1494 = in[335] & in[494];
	wire xformtmp2139;
	assign xformtmp2139 = in[1191] | xformtmp1494;
	wire xformtmp2176;
	assign xformtmp2176 = in[1224] ^ xformtmp2139;
	wire xformtmp2164;
	assign xformtmp2164 = xformtmp1265 & xformtmp2176;
	wire xformtmp1716;
	assign xformtmp1716 = in[781] & xformtmp2164;
	wire xformtmp1916;
	assign xformtmp1916 = in[426] | xformtmp1716;
	wire xformtmp1962;
	assign xformtmp1962 = in[868] | in[904];
	wire xformtmp2021;
	assign xformtmp2021 = xformtmp1916 | xformtmp1962;
	wire xformtmp1460;
	assign xformtmp1460 = in[363] | in[840];
	wire xformtmp1447;
	assign xformtmp1447 = in[1137] & xformtmp1460;
	wire xformtmp2041;
	assign xformtmp2041 = in[271] | in[1102];
	wire xformtmp2214;
	assign xformtmp2214 = in[1129] ^ xformtmp2041;
	wire xformtmp1319;
	assign xformtmp1319 = xformtmp1447 ^ xformtmp2214;
	wire xformtmp1387;
	assign xformtmp1387 = in[1019] ^ in[1145];
	wire xformtmp1620;
	assign xformtmp1620 = xformtmp1319 | xformtmp1387;
	wire xformtmp1846;
	assign xformtmp1846 = in[1424] | xformtmp1620;
	wire xformtmp2238;
	assign xformtmp2238 = in[1251] & xformtmp1846;
	wire xformtmp1313;
	assign xformtmp1313 = xformtmp2021 & xformtmp2238;
	wire xformtmp2003;
	assign xformtmp2003 = in[410] ^ in[789];
	wire xformtmp1297;
	assign xformtmp1297 = in[609] | xformtmp2003;
	wire xformtmp1491;
	assign xformtmp1491 = in[1347] & xformtmp1297;
	wire xformtmp1505;
	assign xformtmp1505 = in[244] | in[398];
	wire xformtmp1760;
	assign xformtmp1760 = in[907] ^ in[1038];
	wire xformtmp1649;
	assign xformtmp1649 = xformtmp1505 & xformtmp1760;
	wire xformtmp1306;
	assign xformtmp1306 = xformtmp1491 & xformtmp1649;
	wire xformtmp1247;
	assign xformtmp1247 = in[394] ^ in[546];
	wire xformtmp1253;
	assign xformtmp1253 = in[312] | in[1252];
	wire xformtmp2050;
	assign xformtmp2050 = in[875] ^ xformtmp1253;
	wire xformtmp1658;
	assign xformtmp1658 = in[278] & xformtmp2050;
	wire xformtmp1528;
	assign xformtmp1528 = in[40] & in[154];
	wire xformtmp2231;
	assign xformtmp2231 = in[873] & xformtmp1528;
	wire xformtmp1884;
	assign xformtmp1884 = in[834] | xformtmp2231;
	wire xformtmp1702;
	assign xformtmp1702 = in[1105] ^ xformtmp1884;
	wire xformtmp2062;
	assign xformtmp2062 = xformtmp1658 | xformtmp1702;
	wire xformtmp2197;
	assign xformtmp2197 = in[1401] | xformtmp2062;
	wire xformtmp2122;
	assign xformtmp2122 = in[58] ^ xformtmp2197;
	wire xformtmp2182;
	assign xformtmp2182 = xformtmp1247 ^ xformtmp2122;
	wire xformtmp1819;
	assign xformtmp1819 = xformtmp1306 ^ xformtmp2182;
	wire xformtmp1511;
	assign xformtmp1511 = xformtmp1313 & xformtmp1819;
	wire xformtmp1654;
	assign xformtmp1654 = in[724] | in[1371];
	wire xformtmp1773;
	assign xformtmp1773 = in[133] | in[139];
	wire xformtmp1973;
	assign xformtmp1973 = in[344] ^ in[1492];
	wire xformtmp1362;
	assign xformtmp1362 = xformtmp1773 ^ xformtmp1973;
	wire xformtmp1478;
	assign xformtmp1478 = in[1096] ^ in[1273];
	wire xformtmp1515;
	assign xformtmp1515 = in[165] & xformtmp1478;
	wire xformtmp1414;
	assign xformtmp1414 = in[229] | in[1208];
	wire xformtmp1707;
	assign xformtmp1707 = in[183] ^ xformtmp1414;
	wire xformtmp2066;
	assign xformtmp2066 = xformtmp1515 | xformtmp1707;
	wire xformtmp1587;
	assign xformtmp1587 = in[827] | in[1324];
	wire xformtmp1748;
	assign xformtmp1748 = in[373] & xformtmp1587;
	wire xformtmp1295;
	assign xformtmp1295 = in[95] | xformtmp1748;
	wire xformtmp1670;
	assign xformtmp1670 = in[831] & in[1153];
	wire xformtmp1849;
	assign xformtmp1849 = xformtmp1295 | xformtmp1670;
	wire xformtmp2241;
	assign xformtmp2241 = in[507] ^ xformtmp1849;
	wire xformtmp1498;
	assign xformtmp1498 = xformtmp2066 & xformtmp2241;
	wire xformtmp1971;
	assign xformtmp1971 = xformtmp1362 ^ xformtmp1498;
	wire xformtmp1762;
	assign xformtmp1762 = in[912] & in[928];
	wire xformtmp1516;
	assign xformtmp1516 = in[631] ^ in[1249];
	wire xformtmp1289;
	assign xformtmp1289 = in[1126] ^ xformtmp1516;
	wire xformtmp1691;
	assign xformtmp1691 = in[51] ^ in[247];
	wire xformtmp2033;
	assign xformtmp2033 = in[127] | in[470];
	wire xformtmp1774;
	assign xformtmp1774 = in[160] ^ xformtmp2033;
	wire xformtmp1966;
	assign xformtmp1966 = xformtmp1691 | xformtmp1774;
	wire xformtmp2020;
	assign xformtmp2020 = in[101] & in[180];
	wire xformtmp1875;
	assign xformtmp1875 = xformtmp1966 ^ xformtmp2020;
	wire xformtmp2208;
	assign xformtmp2208 = xformtmp1289 | xformtmp1875;
	wire xformtmp1379;
	assign xformtmp1379 = xformtmp1762 & xformtmp2208;
	wire xformtmp2018;
	assign xformtmp2018 = in[317] | xformtmp1379;
	wire xformtmp1776;
	assign xformtmp1776 = xformtmp1971 ^ xformtmp2018;
	wire xformtmp1438;
	assign xformtmp1438 = xformtmp1654 | xformtmp1776;
	wire xformtmp1277;
	assign xformtmp1277 = in[797] & in[932];
	wire xformtmp1611;
	assign xformtmp1611 = in[153] & xformtmp1277;
	wire xformtmp1623;
	assign xformtmp1623 = in[389] & in[1256];
	wire xformtmp2245;
	assign xformtmp2245 = in[1297] & xformtmp1623;
	wire xformtmp2159;
	assign xformtmp2159 = in[1000] ^ xformtmp2245;
	wire xformtmp1392;
	assign xformtmp1392 = xformtmp1611 & xformtmp2159;
	wire xformtmp1300;
	assign xformtmp1300 = in[521] | in[765];
	wire xformtmp2004;
	assign xformtmp2004 = in[280] & in[886];
	wire xformtmp1390;
	assign xformtmp1390 = in[1446] | xformtmp2004;
	wire xformtmp1882;
	assign xformtmp1882 = xformtmp1300 ^ xformtmp1390;
	wire xformtmp1370;
	assign xformtmp1370 = in[321] | in[1346];
	wire xformtmp2078;
	assign xformtmp2078 = in[1194] ^ xformtmp1370;
	wire xformtmp2108;
	assign xformtmp2108 = xformtmp1882 | xformtmp2078;
	wire xformtmp1877;
	assign xformtmp1877 = in[331] | xformtmp2108;
	wire xformtmp1530;
	assign xformtmp1530 = xformtmp1392 ^ xformtmp1877;
	wire xformtmp1312;
	assign xformtmp1312 = xformtmp1438 & xformtmp1530;
	wire xformtmp2253;
	assign xformtmp2253 = in[401] & in[661];
	wire xformtmp1864;
	assign xformtmp1864 = in[832] ^ xformtmp2253;
	wire xformtmp1907;
	assign xformtmp1907 = in[814] & xformtmp1864;
	wire xformtmp1720;
	assign xformtmp1720 = in[206] | in[1056];
	wire xformtmp1672;
	assign xformtmp1672 = in[313] & xformtmp1720;
	wire xformtmp1910;
	assign xformtmp1910 = in[196] & in[911];
	wire xformtmp1417;
	assign xformtmp1417 = xformtmp1672 ^ xformtmp1910;
	wire xformtmp2194;
	assign xformtmp2194 = in[288] ^ in[761];
	wire xformtmp1357;
	assign xformtmp1357 = xformtmp1417 ^ xformtmp2194;
	wire xformtmp1775;
	assign xformtmp1775 = in[716] ^ in[850];
	wire xformtmp2011;
	assign xformtmp2011 = xformtmp1357 | xformtmp1775;
	wire xformtmp1468;
	assign xformtmp1468 = xformtmp1907 | xformtmp2011;
	wire xformtmp1999;
	assign xformtmp1999 = in[514] | in[1259];
	wire xformtmp1342;
	assign xformtmp1342 = xformtmp1468 | xformtmp1999;
	wire xformtmp1713;
	assign xformtmp1713 = xformtmp1312 & xformtmp1342;
	wire xformtmp2193;
	assign xformtmp2193 = in[434] ^ in[1463];
	wire xformtmp1924;
	assign xformtmp1924 = in[639] & xformtmp2193;
	wire xformtmp1506;
	assign xformtmp1506 = in[150] ^ in[717];
	wire xformtmp1941;
	assign xformtmp1941 = in[1155] ^ xformtmp1506;
	wire xformtmp2205;
	assign xformtmp2205 = xformtmp1924 | xformtmp1941;
	wire xformtmp2040;
	assign xformtmp2040 = in[729] & xformtmp2205;
	wire xformtmp1351;
	assign xformtmp1351 = in[848] & in[881];
	wire xformtmp1883;
	assign xformtmp1883 = in[1053] & in[1160];
	wire xformtmp1249;
	assign xformtmp1249 = in[906] & in[1263];
	wire xformtmp1432;
	assign xformtmp1432 = in[367] | in[1069];
	wire xformtmp2052;
	assign xformtmp2052 = xformtmp1249 ^ xformtmp1432;
	wire xformtmp1782;
	assign xformtmp1782 = xformtmp1883 | xformtmp2052;
	wire xformtmp1896;
	assign xformtmp1896 = xformtmp1351 ^ xformtmp1782;
	wire xformtmp1996;
	assign xformtmp1996 = in[522] & in[1198];
	wire xformtmp2101;
	assign xformtmp2101 = in[995] | in[1450];
	wire xformtmp1560;
	assign xformtmp1560 = xformtmp1996 & xformtmp2101;
	wire xformtmp2120;
	assign xformtmp2120 = in[445] | xformtmp1560;
	wire xformtmp1959;
	assign xformtmp1959 = in[459] & xformtmp2120;
	wire xformtmp1268;
	assign xformtmp1268 = xformtmp1896 & xformtmp1959;
	wire xformtmp1975;
	assign xformtmp1975 = in[279] ^ in[1136];
	wire xformtmp1594;
	assign xformtmp1594 = in[224] ^ in[1281];
	wire xformtmp2185;
	assign xformtmp2185 = in[114] | xformtmp1594;
	wire xformtmp1383;
	assign xformtmp1383 = in[1386] | xformtmp2185;
	wire xformtmp2013;
	assign xformtmp2013 = in[1384] & xformtmp1383;
	wire xformtmp1257;
	assign xformtmp1257 = xformtmp1975 | xformtmp2013;
	wire xformtmp1831;
	assign xformtmp1831 = in[357] & in[794];
	wire xformtmp1845;
	assign xformtmp1845 = in[1316] & xformtmp1831;
	wire xformtmp1591;
	assign xformtmp1591 = xformtmp1257 ^ xformtmp1845;
	wire xformtmp1700;
	assign xformtmp1700 = xformtmp1268 ^ xformtmp1591;
	wire xformtmp1349;
	assign xformtmp1349 = in[707] ^ xformtmp1700;
	wire xformtmp1435;
	assign xformtmp1435 = in[553] | in[1050];
	wire xformtmp1318;
	assign xformtmp1318 = in[997] | in[1377];
	wire xformtmp1751;
	assign xformtmp1751 = in[231] & in[1372];
	wire xformtmp1834;
	assign xformtmp1834 = in[643] | xformtmp1751;
	wire xformtmp2142;
	assign xformtmp2142 = in[1063] | xformtmp1834;
	wire xformtmp1902;
	assign xformtmp1902 = xformtmp1318 & xformtmp2142;
	wire xformtmp1451;
	assign xformtmp1451 = in[245] & in[1006];
	wire xformtmp2096;
	assign xformtmp2096 = in[1470] ^ xformtmp1451;
	wire xformtmp1854;
	assign xformtmp1854 = xformtmp1902 ^ xformtmp2096;
	wire xformtmp1858;
	assign xformtmp1858 = xformtmp1435 ^ xformtmp1854;
	wire xformtmp1488;
	assign xformtmp1488 = xformtmp1349 & xformtmp1858;
	wire xformtmp1539;
	assign xformtmp1539 = in[342] & in[1183];
	wire xformtmp1696;
	assign xformtmp1696 = in[915] ^ in[988];
	wire xformtmp1440;
	assign xformtmp1440 = in[914] ^ xformtmp1696;
	wire xformtmp2135;
	assign xformtmp2135 = in[776] | in[1454];
	wire xformtmp1798;
	assign xformtmp1798 = xformtmp1440 | xformtmp2135;
	wire xformtmp2207;
	assign xformtmp2207 = xformtmp1539 | xformtmp1798;
	wire xformtmp1309;
	assign xformtmp1309 = in[372] ^ xformtmp2207;
	wire xformtmp1675;
	assign xformtmp1675 = in[4] | in[191];
	wire xformtmp1904;
	assign xformtmp1904 = in[1433] | xformtmp1675;
	wire xformtmp1752;
	assign xformtmp1752 = xformtmp1309 & xformtmp1904;
	wire xformtmp1575;
	assign xformtmp1575 = in[68] ^ in[1186];
	wire xformtmp1559;
	assign xformtmp1559 = in[217] | xformtmp1575;
	wire xformtmp1489;
	assign xformtmp1489 = in[423] | xformtmp1559;
	wire xformtmp2196;
	assign xformtmp2196 = in[265] | xformtmp1489;
	wire xformtmp1629;
	assign xformtmp1629 = xformtmp1752 & xformtmp2196;
	wire xformtmp2104;
	assign xformtmp2104 = xformtmp1488 ^ xformtmp1629;
	wire xformtmp1442;
	assign xformtmp1442 = xformtmp2040 | xformtmp2104;
	wire xformtmp1582;
	assign xformtmp1582 = in[356] | in[1360];
	wire xformtmp1802;
	assign xformtmp1802 = in[1382] & xformtmp1582;
	wire xformtmp1281;
	assign xformtmp1281 = in[1210] & xformtmp1802;
	wire xformtmp1950;
	assign xformtmp1950 = in[370] | in[1045];
	wire xformtmp1969;
	assign xformtmp1969 = in[12] ^ in[1008];
	wire xformtmp1960;
	assign xformtmp1960 = xformtmp1950 ^ xformtmp1969;
	wire xformtmp1655;
	assign xformtmp1655 = in[353] & xformtmp1960;
	wire xformtmp1396;
	assign xformtmp1396 = in[117] ^ xformtmp1655;
	wire xformtmp1757;
	assign xformtmp1757 = in[961] & in[1368];
	wire xformtmp1974;
	assign xformtmp1974 = in[243] & in[1111];
	wire xformtmp1477;
	assign xformtmp1477 = xformtmp1757 & xformtmp1974;
	wire xformtmp2179;
	assign xformtmp2179 = in[1055] ^ in[1304];
	wire xformtmp1788;
	assign xformtmp1788 = in[786] ^ xformtmp2179;
	wire xformtmp1712;
	assign xformtmp1712 = in[1398] | xformtmp1788;
	wire xformtmp2067;
	assign xformtmp2067 = xformtmp1477 & xformtmp1712;
	wire xformtmp1893;
	assign xformtmp1893 = xformtmp1396 & xformtmp2067;
	wire xformtmp2064;
	assign xformtmp2064 = in[186] | in[263];
	wire xformtmp1330;
	assign xformtmp1330 = in[1225] & xformtmp2064;
	wire xformtmp1458;
	assign xformtmp1458 = in[233] ^ in[382];
	wire xformtmp1803;
	assign xformtmp1803 = xformtmp1330 & xformtmp1458;
	wire xformtmp2209;
	assign xformtmp2209 = in[379] | xformtmp1803;
	wire xformtmp2186;
	assign xformtmp2186 = in[454] | xformtmp2209;
	wire xformtmp1301;
	assign xformtmp1301 = xformtmp1893 ^ xformtmp2186;
	wire xformtmp1359;
	assign xformtmp1359 = in[658] & in[993];
	wire xformtmp1285;
	assign xformtmp1285 = in[611] | xformtmp1359;
	wire xformtmp1614;
	assign xformtmp1614 = in[8] ^ in[269];
	wire xformtmp1368;
	assign xformtmp1368 = xformtmp1285 | xformtmp1614;
	wire xformtmp1328;
	assign xformtmp1328 = xformtmp1301 | xformtmp1368;
	wire xformtmp2138;
	assign xformtmp2138 = in[989] ^ in[1397];
	wire xformtmp1870;
	assign xformtmp1870 = in[197] | xformtmp2138;
	wire xformtmp1988;
	assign xformtmp1988 = xformtmp1328 | xformtmp1870;
	wire xformtmp1456;
	assign xformtmp1456 = in[1209] ^ xformtmp1988;
	wire xformtmp1408;
	assign xformtmp1408 = xformtmp1281 | xformtmp1456;
	wire xformtmp1527;
	assign xformtmp1527 = in[728] & in[1052];
	wire xformtmp1943;
	assign xformtmp1943 = in[345] & in[1093];
	wire xformtmp2022;
	assign xformtmp2022 = xformtmp1527 & xformtmp1943;
	wire xformtmp1793;
	assign xformtmp1793 = xformtmp1408 | xformtmp2022;
	wire xformtmp1366;
	assign xformtmp1366 = in[792] | in[1444];
	wire xformtmp1565;
	assign xformtmp1565 = in[607] ^ xformtmp1366;
	wire xformtmp1453;
	assign xformtmp1453 = in[509] & in[978];
	wire xformtmp1680;
	assign xformtmp1680 = in[242] ^ in[1203];
	wire xformtmp2200;
	assign xformtmp2200 = in[1296] & xformtmp1680;
	wire xformtmp1597;
	assign xformtmp1597 = in[795] | in[901];
	wire xformtmp2015;
	assign xformtmp2015 = in[1114] & in[1490];
	wire xformtmp2172;
	assign xformtmp2172 = in[1120] & in[1223];
	wire xformtmp2123;
	assign xformtmp2123 = xformtmp2015 ^ xformtmp2172;
	wire xformtmp2084;
	assign xformtmp2084 = xformtmp1597 ^ xformtmp2123;
	wire xformtmp1284;
	assign xformtmp1284 = in[1192] & xformtmp2084;
	wire xformtmp1504;
	assign xformtmp1504 = in[44] ^ in[376];
	wire xformtmp1709;
	assign xformtmp1709 = in[580] & in[685];
	wire xformtmp2227;
	assign xformtmp2227 = xformtmp1504 | xformtmp1709;
	wire xformtmp1703;
	assign xformtmp1703 = in[334] | xformtmp2227;
	wire xformtmp1409;
	assign xformtmp1409 = xformtmp1284 ^ xformtmp1703;
	wire xformtmp1953;
	assign xformtmp1953 = in[615] | in[1211];
	wire xformtmp1278;
	assign xformtmp1278 = in[1140] & xformtmp1953;
	wire xformtmp1865;
	assign xformtmp1865 = in[466] | in[1015];
	wire xformtmp2088;
	assign xformtmp2088 = xformtmp1278 | xformtmp1865;
	wire xformtmp2228;
	assign xformtmp2228 = xformtmp1409 ^ xformtmp2088;
	wire xformtmp1425;
	assign xformtmp1425 = xformtmp2200 & xformtmp2228;
	wire xformtmp2255;
	assign xformtmp2255 = in[764] | xformtmp1425;
	wire xformtmp1711;
	assign xformtmp1711 = xformtmp1453 ^ xformtmp2255;
	wire xformtmp1612;
	assign xformtmp1612 = in[104] | in[686];
	wire xformtmp1721;
	assign xformtmp1721 = in[576] ^ in[1467];
	wire xformtmp1619;
	assign xformtmp1619 = in[1170] & xformtmp1721;
	wire xformtmp1800;
	assign xformtmp1800 = xformtmp1612 ^ xformtmp1619;
	wire xformtmp1928;
	assign xformtmp1928 = in[1030] ^ in[1270];
	wire xformtmp2117;
	assign xformtmp2117 = xformtmp1800 ^ xformtmp1928;
	wire xformtmp1624;
	assign xformtmp1624 = xformtmp1711 ^ xformtmp2117;
	wire xformtmp2147;
	assign xformtmp2147 = xformtmp1565 & xformtmp1624;
	wire xformtmp1270;
	assign xformtmp1270 = xformtmp1793 ^ xformtmp2147;
	wire xformtmp1524;
	assign xformtmp1524 = in[677] & in[1103];
	wire xformtmp1684;
	assign xformtmp1684 = in[391] & xformtmp1524;
	wire xformtmp1507;
	assign xformtmp1507 = in[214] & xformtmp1684;
	wire xformtmp1446;
	assign xformtmp1446 = in[31] | xformtmp1507;
	wire xformtmp1422;
	assign xformtmp1422 = in[900] & xformtmp1446;
	wire xformtmp1294;
	assign xformtmp1294 = xformtmp1270 ^ xformtmp1422;
	wire xformtmp1967;
	assign xformtmp1967 = in[869] | in[1238];
	wire xformtmp1554;
	assign xformtmp1554 = in[326] & xformtmp1967;
	wire xformtmp1947;
	assign xformtmp1947 = in[1193] | in[1355];
	wire xformtmp1683;
	assign xformtmp1683 = in[1351] ^ xformtmp1947;
	wire xformtmp1897;
	assign xformtmp1897 = xformtmp1554 & xformtmp1683;
	wire xformtmp1305;
	assign xformtmp1305 = in[171] | in[768];
	wire xformtmp1818;
	assign xformtmp1818 = in[956] ^ xformtmp1305;
	wire xformtmp1323;
	assign xformtmp1323 = in[877] ^ in[990];
	wire xformtmp1452;
	assign xformtmp1452 = in[482] | xformtmp1323;
	wire xformtmp2222;
	assign xformtmp2222 = in[1132] & xformtmp1452;
	wire xformtmp1906;
	assign xformtmp1906 = xformtmp1818 & xformtmp2222;
	wire xformtmp1492;
	assign xformtmp1492 = xformtmp1897 & xformtmp1906;
	wire xformtmp1476;
	assign xformtmp1476 = in[177] | in[760];
	wire xformtmp1698;
	assign xformtmp1698 = in[223] ^ xformtmp1476;
	wire xformtmp1770;
	assign xformtmp1770 = in[706] | xformtmp1698;
	wire xformtmp2247;
	assign xformtmp2247 = in[239] & in[1081];
	wire xformtmp1393;
	assign xformtmp1393 = xformtmp1770 | xformtmp2247;
	wire xformtmp1961;
	assign xformtmp1961 = in[718] | xformtmp1393;
	wire xformtmp1598;
	assign xformtmp1598 = xformtmp1492 & xformtmp1961;
	wire xformtmp1445;
	assign xformtmp1445 = xformtmp1294 | xformtmp1598;
	wire xformtmp2252;
	assign xformtmp2252 = xformtmp1442 | xformtmp1445;
	wire xformtmp2001;
	assign xformtmp2001 = xformtmp1713 & xformtmp2252;
	wire xformtmp1663;
	assign xformtmp1663 = xformtmp1511 | xformtmp2001;
	assign out[499] = xformtmp1391 & xformtmp1663;
endmodule

module tb();
    reg[499:0] results[1];
    reg[1499:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%1500b]", data[0]);
        #1
        $display("results = [%500b]", results[0]);
        $writememb("results.txt", results);
    end
endmodule

