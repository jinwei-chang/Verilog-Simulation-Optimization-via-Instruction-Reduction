module dut (out, in);
	output[6:0] out;
	input[35:0] in;
	wire origtmp1;
	wire origtmp2;
	wire origtmp3;
	wire origtmp4;
	wire origtmp5;
	wire origtmp6;
	wire origtmp7;
	wire origtmp8;
	wire origtmp9;
	wire origtmp10;
	wire origtmp11;
	wire origtmp12;
	wire origtmp13;
	wire origtmp14;
	wire origtmp15;
	wire origtmp16;
	wire origtmp17;
	wire origtmp18;
	wire origtmp19;
	wire origtmp20;
	wire origtmp21;
	wire origtmp22;
	wire origtmp23;
	wire origtmp24;
	wire origtmp25;
	wire origtmp26;
	wire origtmp27;
	wire origtmp28;
	wire origtmp29;
	wire origtmp30;
	wire origtmp31;
	wire origtmp32;
	wire origtmp33;
	wire origtmp34;
	wire origtmp35;
	wire origtmp36;
	wire origtmp37;
	wire origtmp38;
	wire origtmp39;
	wire origtmp40;
	wire origtmp41;
	wire origtmp42;
	wire origtmp43;
	wire origtmp44;
	wire origtmp45;
	wire origtmp46;
	wire origtmp47;
	wire origtmp48;
	wire origtmp49;
	wire origtmp50;
	wire origtmp51;
	wire origtmp52;
	wire origtmp53;
	wire origtmp54;
	wire origtmp55;
	wire origtmp56;
	wire origtmp57;
	wire origtmp58;
	wire origtmp59;
	wire origtmp60;
	wire origtmp61;
	wire origtmp62;
	wire origtmp63;
	wire origtmp64;
	wire origtmp65;
	wire origtmp66;
	wire origtmp67;
	wire origtmp68;
	wire origtmp69;
	wire origtmp70;
	wire origtmp71;
	wire origtmp72;
	wire origtmp73;
	wire origtmp74;
	wire origtmp75;
	wire origtmp76;
	wire origtmp77;
	wire origtmp78;
	wire origtmp79;
	wire origtmp80;
	wire origtmp81;
	wire origtmp82;
	wire origtmp83;
	wire origtmp84;
	wire origtmp85;
	wire origtmp86;
	wire origtmp87;
	wire origtmp88;
	wire origtmp89;
	wire origtmp90;
	wire origtmp91;
	wire origtmp92;
	wire origtmp93;
	wire origtmp94;
	wire origtmp95;
	wire origtmp96;
	wire origtmp97;
	wire origtmp98;
	wire origtmp99;
	wire origtmp100;
	wire origtmp101;
	wire origtmp102;
	wire origtmp103;
	wire origtmp104;
	wire origtmp105;
	wire origtmp106;
	wire origtmp107;
	wire origtmp108;
	wire origtmp109;
	wire origtmp110;
	wire origtmp111;
	wire origtmp112;
	wire origtmp113;
	wire origtmp114;
	wire origtmp115;
	wire origtmp116;
	wire origtmp117;
	wire origtmp118;
	wire origtmp119;
	wire origtmp120;
	wire origtmp121;
	wire origtmp122;
	wire origtmp123;
	wire origtmp124;
	wire origtmp125;
	wire origtmp126;
	wire origtmp127;
	wire origtmp128;
	wire origtmp129;
	wire origtmp130;
	wire origtmp131;
	wire origtmp132;
	wire origtmp133;
	wire origtmp134;
	wire origtmp135;
	wire origtmp136;
	wire origtmp137;
	wire origtmp138;
	wire origtmp139;
	wire origtmp140;
	wire origtmp141;
	wire origtmp142;
	wire origtmp143;
	wire origtmp144;
	wire origtmp145;
	wire origtmp146;
	wire origtmp147;
	wire origtmp148;
	wire origtmp149;
	wire origtmp150;
	wire origtmp151;
	wire origtmp152;
	wire origtmp153;
	wire origtmp154;
	wire origtmp155;
	wire origtmp156;
	wire origtmp157;
	wire origtmp158;
	wire origtmp159;
	wire origtmp160;
	wire origtmp161;
	wire origtmp162;
	wire origtmp163;
	wire origtmp164;
	wire origtmp165;
	wire origtmp166;
	wire origtmp167;
	wire origtmp168;
	wire origtmp169;
	wire origtmp170;
	wire origtmp171;
	wire origtmp172;
	wire origtmp173;
	wire origtmp174;
	wire origtmp175;
	wire origtmp176;
	wire origtmp177;
	wire origtmp178;
	wire origtmp179;
	wire origtmp180;
	wire origtmp181;
	wire origtmp182;
	wire origtmp183;
	wire origtmp184;
	wire origtmp185;
	wire origtmp186;
	wire origtmp187;
	wire origtmp188;
	wire origtmp189;
	wire origtmp190;
	wire origtmp191;
	wire origtmp192;
	wire origtmp193;
	wire origtmp194;
	wire origtmp195;
	wire origtmp196;
	wire origtmp197;
	wire origtmp198;
	wire origtmp199;
	wire origtmp200;
	wire origtmp201;
	wire origtmp202;
	wire origtmp203;
	wire origtmp204;
	wire origtmp205;
	wire origtmp206;
	wire origtmp207;
	wire origtmp208;
	wire origtmp209;
	wire origtmp210;
	wire origtmp211;
	wire origtmp212;
	wire origtmp213;
	wire origtmp214;
	wire origtmp215;
	wire origtmp216;
	wire origtmp217;
	wire origtmp218;
	wire origtmp219;
	wire origtmp220;
	wire origtmp221;
	wire origtmp222;
	wire origtmp223;
	wire origtmp224;
	wire origtmp225;
	wire origtmp226;
	wire origtmp227;
	wire origtmp228;
	wire origtmp229;
	wire origtmp230;
	wire origtmp231;
	wire origtmp232;
	wire origtmp233;
	wire origtmp234;
	wire origtmp235;
	wire origtmp236;
	wire origtmp237;
	wire origtmp238;
	wire origtmp239;
	wire origtmp240;
	wire origtmp241;
	wire origtmp242;
	wire origtmp243;
	wire origtmp244;
	wire origtmp245;
	wire origtmp246;
	wire origtmp247;
	wire origtmp248;
	wire origtmp249;
	wire origtmp250;
	wire origtmp251;
	wire origtmp252;
	wire origtmp253;
	wire origtmp254;
	wire origtmp255;
	wire origtmp256;
	wire origtmp257;
	wire origtmp258;
	wire origtmp259;
	wire origtmp260;
	wire origtmp261;
	wire origtmp262;
	wire origtmp263;
	wire origtmp264;
	wire origtmp265;
	wire origtmp266;
	wire origtmp267;
	wire origtmp268;
	wire origtmp269;
	wire origtmp270;
	wire origtmp271;
	wire origtmp272;
	wire origtmp273;
	wire origtmp274;
	wire origtmp275;
	wire origtmp276;
	wire origtmp277;
	wire origtmp278;
	wire origtmp279;
	wire origtmp280;
	wire origtmp281;
	wire origtmp282;
	wire origtmp283;
	wire origtmp284;
	wire origtmp285;
	wire origtmp286;
	wire origtmp287;
	wire origtmp288;
	wire origtmp289;
	wire origtmp290;
	wire origtmp291;
	wire origtmp292;
	wire origtmp293;
	wire origtmp294;
	wire origtmp295;
	wire origtmp296;
	wire origtmp297;
	wire origtmp298;
	wire origtmp299;
	wire origtmp300;
	wire origtmp301;
	wire origtmp302;
	wire origtmp303;
	wire origtmp304;
	wire origtmp305;
	wire origtmp306;
	wire origtmp307;
	assign origtmp1 = ~in[0];
	assign origtmp2 = ~in[1];
	assign origtmp3 = ~in[3];
	assign origtmp4 = ~in[5];
	assign origtmp5 = ~in[7];
	assign origtmp6 = ~in[9];
	assign origtmp7 = ~in[11];
	assign origtmp8 = ~in[13];
	assign origtmp9 = ~in[15];
	assign origtmp10 = ~in[17];
	assign origtmp11 = ~in[19];
	assign origtmp12 = ~in[21];
	assign origtmp13 = ~in[23];
	assign origtmp14 = ~in[25];
	assign origtmp15 = ~in[27];
	assign origtmp16 = ~in[29];
	assign origtmp17 = ~in[31];
	assign origtmp18 = ~in[33];
	assign origtmp20 = origtmp1 & in[1];
	assign origtmp19 = ~origtmp20;
	assign origtmp22 = in[2] | origtmp2;
	assign origtmp21 = ~origtmp22;
	assign origtmp24 = in[4] | origtmp2;
	assign origtmp23 = ~origtmp24;
	assign origtmp26 = origtmp3 & in[5];
	assign origtmp25 = ~origtmp26;
	assign origtmp28 = origtmp5 & in[9];
	assign origtmp27 = ~origtmp28;
	assign origtmp30 = origtmp7 & in[13];
	assign origtmp29 = ~origtmp30;
	assign origtmp32 = origtmp9 & in[17];
	assign origtmp31 = ~origtmp32;
	assign origtmp34 = origtmp11 & in[21];
	assign origtmp33 = ~origtmp34;
	assign origtmp36 = origtmp13 & in[25];
	assign origtmp35 = ~origtmp36;
	assign origtmp38 = origtmp15 & in[29];
	assign origtmp37 = ~origtmp38;
	assign origtmp40 = origtmp17 & in[33];
	assign origtmp39 = ~origtmp40;
	assign origtmp42 = in[6] | origtmp4;
	assign origtmp41 = ~origtmp42;
	assign origtmp44 = in[8] | origtmp4;
	assign origtmp43 = ~origtmp44;
	assign origtmp46 = in[10] | origtmp6;
	assign origtmp45 = ~origtmp46;
	assign origtmp48 = in[12] | origtmp6;
	assign origtmp47 = ~origtmp48;
	assign origtmp50 = in[14] | origtmp8;
	assign origtmp49 = ~origtmp50;
	assign origtmp52 = in[16] | origtmp8;
	assign origtmp51 = ~origtmp52;
	assign origtmp54 = in[18] | origtmp10;
	assign origtmp53 = ~origtmp54;
	assign origtmp56 = in[20] | origtmp10;
	assign origtmp55 = ~origtmp56;
	assign origtmp58 = in[22] | origtmp12;
	assign origtmp57 = ~origtmp58;
	assign origtmp60 = in[24] | origtmp12;
	assign origtmp59 = ~origtmp60;
	assign origtmp62 = in[26] | origtmp14;
	assign origtmp61 = ~origtmp62;
	assign origtmp64 = in[28] | origtmp14;
	assign origtmp63 = ~origtmp64;
	assign origtmp66 = in[30] | origtmp16;
	assign origtmp65 = ~origtmp66;
	assign origtmp68 = in[32] | origtmp16;
	assign origtmp67 = ~origtmp68;
	assign origtmp70 = in[34] | origtmp18;
	assign origtmp69 = ~origtmp70;
	assign origtmp72 = in[35] | origtmp18;
	assign origtmp71 = ~origtmp72;
	assign origtmp74 = origtmp37 & origtmp39;
	assign origtmp75 = origtmp74 & origtmp35;
	assign origtmp76 = origtmp75 & origtmp33;
	assign origtmp77 = origtmp76 & origtmp31;
	assign origtmp78 = origtmp77 & origtmp29;
	assign origtmp79 = origtmp78 & origtmp27;
	assign origtmp80 = origtmp79 & origtmp25;
	assign origtmp73 = origtmp80 & origtmp19;
	assign origtmp81 = ~origtmp73;
	assign origtmp82 = ~origtmp73;
	assign out[0] = ~origtmp73;
	assign origtmp83 = origtmp81 ^ origtmp19;
	assign origtmp84 = origtmp81 ^ origtmp25;
	assign origtmp85 = origtmp81 ^ origtmp27;
	assign origtmp86 = origtmp81 ^ origtmp29;
	assign origtmp87 = origtmp81 ^ origtmp31;
	assign origtmp88 = origtmp81 ^ origtmp33;
	assign origtmp90 = in[0] & origtmp82;
	assign origtmp89 = ~origtmp90;
	assign origtmp91 = origtmp81 ^ origtmp35;
	assign origtmp93 = origtmp82 & in[3];
	assign origtmp92 = ~origtmp93;
	assign origtmp94 = origtmp81 ^ origtmp37;
	assign origtmp96 = origtmp82 & in[7];
	assign origtmp95 = ~origtmp96;
	assign origtmp97 = origtmp81 ^ origtmp39;
	assign origtmp99 = origtmp82 & in[11];
	assign origtmp98 = ~origtmp99;
	assign origtmp101 = origtmp82 & in[15];
	assign origtmp100 = ~origtmp101;
	assign origtmp103 = origtmp82 & in[19];
	assign origtmp102 = ~origtmp103;
	assign origtmp105 = origtmp82 & in[23];
	assign origtmp104 = ~origtmp105;
	assign origtmp107 = origtmp82 & in[27];
	assign origtmp106 = ~origtmp107;
	assign origtmp109 = origtmp82 & in[31];
	assign origtmp108 = ~origtmp109;
	assign origtmp111 = origtmp83 & origtmp21;
	assign origtmp110 = ~origtmp111;
	assign origtmp113 = origtmp83 & origtmp23;
	assign origtmp112 = ~origtmp113;
	assign origtmp115 = origtmp84 & origtmp41;
	assign origtmp114 = ~origtmp115;
	assign origtmp117 = origtmp85 & origtmp45;
	assign origtmp116 = ~origtmp117;
	assign origtmp119 = origtmp86 & origtmp49;
	assign origtmp118 = ~origtmp119;
	assign origtmp121 = origtmp87 & origtmp53;
	assign origtmp120 = ~origtmp121;
	assign origtmp123 = origtmp88 & origtmp57;
	assign origtmp122 = ~origtmp123;
	assign origtmp125 = origtmp91 & origtmp61;
	assign origtmp124 = ~origtmp125;
	assign origtmp127 = origtmp94 & origtmp65;
	assign origtmp126 = ~origtmp127;
	assign origtmp129 = origtmp97 & origtmp69;
	assign origtmp128 = ~origtmp129;
	assign origtmp131 = origtmp84 & origtmp43;
	assign origtmp130 = ~origtmp131;
	assign origtmp133 = origtmp85 & origtmp47;
	assign origtmp132 = ~origtmp133;
	assign origtmp135 = origtmp86 & origtmp51;
	assign origtmp134 = ~origtmp135;
	assign origtmp137 = origtmp87 & origtmp55;
	assign origtmp136 = ~origtmp137;
	assign origtmp139 = origtmp88 & origtmp59;
	assign origtmp138 = ~origtmp139;
	assign origtmp141 = origtmp91 & origtmp63;
	assign origtmp140 = ~origtmp141;
	assign origtmp143 = origtmp94 & origtmp67;
	assign origtmp142 = ~origtmp143;
	assign origtmp145 = origtmp97 & origtmp71;
	assign origtmp144 = ~origtmp145;
	assign origtmp147 = origtmp126 & origtmp128;
	assign origtmp148 = origtmp147 & origtmp124;
	assign origtmp149 = origtmp148 & origtmp122;
	assign origtmp150 = origtmp149 & origtmp120;
	assign origtmp151 = origtmp150 & origtmp118;
	assign origtmp152 = origtmp151 & origtmp116;
	assign origtmp153 = origtmp152 & origtmp114;
	assign origtmp146 = origtmp153 & origtmp110;
	assign origtmp154 = ~origtmp112;
	assign origtmp155 = ~origtmp130;
	assign origtmp156 = ~origtmp132;
	assign origtmp157 = ~origtmp134;
	assign origtmp158 = ~origtmp136;
	assign origtmp159 = ~origtmp138;
	assign origtmp160 = ~origtmp140;
	assign origtmp161 = ~origtmp142;
	assign origtmp162 = ~origtmp144;
	assign origtmp163 = ~origtmp146;
	assign origtmp164 = ~origtmp146;
	assign out[1] = ~origtmp146;
	assign origtmp165 = origtmp163 ^ origtmp110;
	assign origtmp166 = origtmp163 ^ origtmp114;
	assign origtmp167 = origtmp163 ^ origtmp116;
	assign origtmp168 = origtmp163 ^ origtmp118;
	assign origtmp170 = in[2] & origtmp164;
	assign origtmp169 = ~origtmp170;
	assign origtmp171 = origtmp163 ^ origtmp120;
	assign origtmp173 = origtmp164 & in[6];
	assign origtmp172 = ~origtmp173;
	assign origtmp174 = origtmp163 ^ origtmp122;
	assign origtmp176 = origtmp164 & in[10];
	assign origtmp175 = ~origtmp176;
	assign origtmp177 = origtmp163 ^ origtmp124;
	assign origtmp179 = origtmp164 & in[14];
	assign origtmp178 = ~origtmp179;
	assign origtmp180 = origtmp163 ^ origtmp126;
	assign origtmp182 = origtmp164 & in[18];
	assign origtmp181 = ~origtmp182;
	assign origtmp183 = origtmp163 ^ origtmp128;
	assign origtmp185 = origtmp164 & in[22];
	assign origtmp184 = ~origtmp185;
	assign origtmp187 = origtmp164 & in[26];
	assign origtmp186 = ~origtmp187;
	assign origtmp189 = origtmp164 & in[30];
	assign origtmp188 = ~origtmp189;
	assign origtmp191 = origtmp164 & in[34];
	assign origtmp190 = ~origtmp191;
	assign origtmp193 = origtmp165 & origtmp154;
	assign origtmp192 = ~origtmp193;
	assign origtmp195 = origtmp166 & origtmp155;
	assign origtmp194 = ~origtmp195;
	assign origtmp197 = origtmp167 & origtmp156;
	assign origtmp196 = ~origtmp197;
	assign origtmp199 = origtmp168 & origtmp157;
	assign origtmp198 = ~origtmp199;
	assign origtmp201 = origtmp171 & origtmp158;
	assign origtmp200 = ~origtmp201;
	assign origtmp203 = origtmp174 & origtmp159;
	assign origtmp202 = ~origtmp203;
	assign origtmp205 = origtmp177 & origtmp160;
	assign origtmp204 = ~origtmp205;
	assign origtmp207 = origtmp180 & origtmp161;
	assign origtmp206 = ~origtmp207;
	assign origtmp209 = origtmp183 & origtmp162;
	assign origtmp208 = ~origtmp209;
	assign origtmp211 = origtmp206 & origtmp208;
	assign origtmp212 = origtmp211 & origtmp204;
	assign origtmp213 = origtmp212 & origtmp202;
	assign origtmp214 = origtmp213 & origtmp200;
	assign origtmp215 = origtmp214 & origtmp198;
	assign origtmp216 = origtmp215 & origtmp196;
	assign origtmp217 = origtmp216 & origtmp194;
	assign origtmp210 = origtmp217 & origtmp192;
	assign origtmp218 = ~origtmp210;
	assign out[2] = ~origtmp210;
	assign origtmp220 = in[4] & origtmp218;
	assign origtmp219 = ~origtmp220;
	assign origtmp222 = origtmp218 & in[8];
	assign origtmp221 = ~origtmp222;
	assign origtmp224 = origtmp218 & in[12];
	assign origtmp223 = ~origtmp224;
	assign origtmp226 = origtmp218 & in[16];
	assign origtmp225 = ~origtmp226;
	assign origtmp228 = origtmp218 & in[20];
	assign origtmp227 = ~origtmp228;
	assign origtmp230 = origtmp218 & in[24];
	assign origtmp229 = ~origtmp230;
	assign origtmp232 = origtmp218 & in[28];
	assign origtmp231 = ~origtmp232;
	assign origtmp234 = origtmp218 & in[32];
	assign origtmp233 = ~origtmp234;
	assign origtmp236 = origtmp218 & in[35];
	assign origtmp235 = ~origtmp236;
	assign origtmp238 = origtmp169 & origtmp219;
	assign origtmp239 = origtmp238 & origtmp89;
	assign origtmp240 = origtmp239 & in[1];
	assign origtmp237 = ~origtmp240;
	assign origtmp242 = origtmp221 & in[5];
	assign origtmp243 = origtmp242 & origtmp172;
	assign origtmp244 = origtmp243 & origtmp92;
	assign origtmp241 = ~origtmp244;
	assign origtmp246 = origtmp223 & in[9];
	assign origtmp247 = origtmp246 & origtmp175;
	assign origtmp248 = origtmp247 & origtmp95;
	assign origtmp245 = ~origtmp248;
	assign origtmp250 = origtmp225 & in[13];
	assign origtmp251 = origtmp250 & origtmp178;
	assign origtmp252 = origtmp251 & origtmp98;
	assign origtmp249 = ~origtmp252;
	assign origtmp254 = origtmp227 & in[17];
	assign origtmp255 = origtmp254 & origtmp181;
	assign origtmp256 = origtmp255 & origtmp100;
	assign origtmp253 = ~origtmp256;
	assign origtmp258 = origtmp229 & in[21];
	assign origtmp259 = origtmp258 & origtmp184;
	assign origtmp260 = origtmp259 & origtmp102;
	assign origtmp257 = ~origtmp260;
	assign origtmp262 = origtmp231 & in[25];
	assign origtmp263 = origtmp262 & origtmp186;
	assign origtmp264 = origtmp263 & origtmp104;
	assign origtmp261 = ~origtmp264;
	assign origtmp266 = origtmp233 & in[29];
	assign origtmp267 = origtmp266 & origtmp188;
	assign origtmp268 = origtmp267 & origtmp106;
	assign origtmp265 = ~origtmp268;
	assign origtmp270 = origtmp235 & in[33];
	assign origtmp271 = origtmp270 & origtmp190;
	assign origtmp272 = origtmp271 & origtmp108;
	assign origtmp269 = ~origtmp272;
	assign origtmp273 = ~origtmp237;
	assign origtmp275 = origtmp265 & origtmp269;
	assign origtmp276 = origtmp275 & origtmp261;
	assign origtmp277 = origtmp276 & origtmp257;
	assign origtmp278 = origtmp277 & origtmp253;
	assign origtmp279 = origtmp278 & origtmp249;
	assign origtmp280 = origtmp279 & origtmp245;
	assign origtmp274 = origtmp280 & origtmp241;
	assign origtmp281 = ~origtmp249;
	assign origtmp282 = ~origtmp257;
	assign origtmp283 = ~origtmp261;
	assign origtmp284 = ~origtmp265;
	assign origtmp285 = origtmp273 | origtmp274;
	assign out[3] = ~origtmp285;
	assign origtmp287 = origtmp245 & origtmp281;
	assign origtmp286 = ~origtmp287;
	assign origtmp289 = origtmp282 & origtmp253;
	assign origtmp290 = origtmp289 & origtmp249;
	assign origtmp291 = origtmp290 & origtmp245;
	assign origtmp288 = ~origtmp291;
	assign origtmp293 = origtmp249 & origtmp283;
	assign origtmp294 = origtmp293 & origtmp253;
	assign origtmp292 = ~origtmp294;
	assign origtmp296 = origtmp261 & origtmp284;
	assign origtmp297 = origtmp296 & origtmp249;
	assign origtmp298 = origtmp297 & origtmp245;
	assign origtmp295 = ~origtmp298;
	assign origtmp299 = origtmp286 & origtmp253;
	assign origtmp300 = origtmp299 & origtmp245;
	assign origtmp301 = origtmp300 & origtmp241;
	assign out[4] = ~origtmp301;
	assign origtmp302 = origtmp288 & origtmp292;
	assign origtmp303 = origtmp302 & origtmp245;
	assign origtmp304 = origtmp303 & origtmp241;
	assign out[5] = ~origtmp304;
	assign origtmp305 = origtmp288 & origtmp295;
	assign origtmp306 = origtmp305 & origtmp286;
	assign origtmp307 = origtmp306 & origtmp241;
	assign out[6] = ~origtmp307;
endmodule

module tb();
    reg[6:0] results[1];
    reg[35:0] data[1];
    dut duttest(results[0], data[0]);
    initial begin
        $readmemb("data.txt", data);
        $display("data = [%36b]", data[0]);
        #1
        $display("results = [%7b]", results[0]);
        $writememb("results.txt", results);
    end
endmodule

